

real kernel_1_re[4][1][3][3] =
    '{'{'{  '{0.1539, 0.1462, 0.1500},
            '{0.1833, 0.1852, 0.1734},
            '{0.1660, 0.1688, 0.1406}}},
        '{'{'{0.1565, 0.1589, 0.1283},
            '{0.1880, 0.2126, 0.1786},
            '{0.1511, 0.1563, 0.1618}}},
        '{'{'{0.1212, 0.1438, 0.1486},
            '{0.1760, 0.1886, 0.1718},
            '{0.1556, 0.1773, 0.1559}}},
        '{'{'{0.1446, 0.1665, 0.1416},
            '{0.1583, 0.1853, 0.1838},
            '{0.1626, 0.1682, 0.1605}}}};

real conv_1_bias_re[4] = '{0.0042, 0.0091, 0.0215, 0.0043};

real kernel_2_re[8][4][3][3] =
'{'{'{'{-0.0319, -0.1899, -0.2296},
          '{ 0.1554,  0.0842,  0.0591},
          '{ 0.1143,  0.1015,  0.1385}},

         '{'{-0.0157, -0.1726, -0.2313},
          '{ 0.1664,  0.0872,  0.0769},
          '{ 0.1083,  0.1119,  0.1464}},

         '{'{ 0.0011, -0.1682, -0.2138},
          '{ 0.1637,  0.0784,  0.1035},
          '{ 0.1004,  0.1030,  0.1469}},

         '{'{-0.0148, -0.1645, -0.2315},
          '{ 0.1349,  0.0929,  0.0954},
          '{ 0.1055,  0.1180,  0.1644}}},


        '{'{'{ 0.1411,  0.1692,  0.1972},
          '{-0.0381, -0.0073, -0.0471},
          '{-0.2295, -0.2062, -0.1685}},

         '{'{ 0.1446,  0.1645,  0.2036},
          '{-0.0178, -0.0142, -0.0356},
          '{-0.2265, -0.2035, -0.1789}},

         '{'{ 0.1558,  0.1740,  0.1710},
          '{-0.0281,  0.0020, -0.0508},
          '{-0.2131, -0.1881, -0.1271}},

         '{'{ 0.1296,  0.1759,  0.1908},
          '{-0.0244, -0.0053, -0.0315},
          '{-0.2371, -0.2070, -0.1888}}},


        '{'{'{ 0.1123,  0.1737,  0.1293},
          '{-0.1358, -0.0241,  0.1197},
          '{-0.1039, -0.0048,  0.1370}},

         '{'{ 0.1034,  0.1656,  0.1651},
          '{-0.1422, -0.0308,  0.1236},
          '{-0.0973, -0.0021,  0.1276}},

         '{'{ 0.1150,  0.1635,  0.1397},
          '{-0.0980, -0.0120,  0.1381},
          '{-0.1031,  0.0399,  0.1589}},

         '{'{ 0.1170,  0.1584,  0.1422},
          '{-0.1272, -0.0166,  0.1201},
          '{-0.0965, -0.0030,  0.1398}}},


        '{'{'{-0.2190, -0.0268,  0.1735},
          '{-0.2396,  0.0768,  0.1452},
          '{-0.0890,  0.1065,  0.1142}},

         '{'{-0.2326, -0.0030,  0.1862},
          '{-0.2336,  0.1006,  0.1250},
          '{-0.1130,  0.0963,  0.0891}},

         '{'{-0.2285, -0.0143,  0.1712},
          '{-0.2385,  0.0702,  0.1299},
          '{-0.1003,  0.1191,  0.0898}},

         '{'{-0.2438, -0.0075,  0.1883},
          '{-0.2146,  0.0926,  0.1272},
          '{-0.0989,  0.1199,  0.0957}}},


        '{'{'{ 0.0889,  0.0774,  0.0695},
          '{ 0.0789,  0.0695,  0.0272},
          '{ 0.0723,  0.0601,  0.0774}},

         '{'{ 0.0776,  0.0805,  0.1091},
          '{ 0.0525,  0.0440,  0.0401},
          '{ 0.0810,  0.0173,  0.0697}},

         '{'{ 0.0998,  0.1011,  0.0751},
          '{ 0.0580,  0.0490,  0.0298},
          '{ 0.0617,  0.0381,  0.0560}},

         '{'{ 0.0821,  0.0954,  0.0745},
          '{ 0.0504,  0.0512,  0.0298},
          '{ 0.0640,  0.0590,  0.0566}}},


        '{'{'{ 0.0847,  0.0913,  0.0957},
          '{ 0.0715,  0.1075,  0.1650},
          '{-0.2236, -0.2098, -0.0789}},

         '{'{ 0.1168,  0.0894,  0.1131},
          '{ 0.0702,  0.1093,  0.1502},
          '{-0.2244, -0.2079, -0.0612}},

         '{'{ 0.1050,  0.0908,  0.1138},
          '{ 0.0856,  0.0972,  0.1717},
          '{-0.2092, -0.2137, -0.0616}},

         '{'{ 0.1140,  0.0951,  0.0960},
          '{ 0.0552,  0.1049,  0.1738},
          '{-0.2246, -0.2185, -0.0448}}},


        '{'{'{-0.0724,  0.0585,  0.1229},
          '{ 0.1074,  0.0943,  0.0977},
          '{ 0.1079,  0.0679,  0.0185}},

         '{'{-0.0698,  0.0369,  0.1319},
          '{ 0.1020,  0.0863,  0.0851},
          '{ 0.1065,  0.0726, -0.0036}},

         '{'{-0.0626,  0.0799,  0.1400},
          '{ 0.1335,  0.1000,  0.0918},
          '{ 0.1321,  0.0766, -0.0242}},

         '{'{-0.0550,  0.0739,  0.1409},
          '{ 0.1115,  0.0998,  0.0818},
          '{ 0.1072,  0.0528, -0.0006}}},


        '{'{'{ 0.0384,  0.0845,  0.0903},
          '{ 0.0639,  0.0779,  0.0469},
          '{ 0.0918,  0.0794,  0.0989}},

         '{'{ 0.0329,  0.0884,  0.1046},
          '{ 0.0715,  0.0581,  0.0796},
          '{ 0.0852,  0.0732,  0.0875}},

         '{'{ 0.0617,  0.0848,  0.0762},
          '{ 0.0824,  0.0857,  0.0346},
          '{ 0.0783,  0.0761,  0.0680}},

         '{'{ 0.0630,  0.0906,  0.1090},
          '{ 0.0751,  0.0786,  0.0512},
          '{ 0.0778,  0.0762,  0.0936}}}};


real conv_2_bias_re[8] = '{ 0.0133,  0.0802,  0.0038, -0.0109,  0.0106,  0.0513, -0.0028,  0.0026};

real fc1_weights_re[64][200] = '{'{ 1.4964e-02,  1.6226e-01, -9.3647e-03, -1.8295e-02, -2.4734e-03,
         -1.8522e-02, -9.0810e-02, -1.8042e-01, -1.5219e-01, -5.3419e-02,
         -3.2822e-02,  8.5469e-02,  1.8318e-01,  4.7955e-02,  8.1632e-02,
         -1.5248e-02,  1.5170e-01,  1.3182e-01,  6.6886e-02, -1.0131e-01,
         -1.4351e-01,  1.2600e-03,  5.3629e-02,  8.9052e-02, -2.0993e-02,
         -1.1332e-01,  1.5099e-02, -1.8489e-02,  2.6553e-02, -1.9306e-01,
         -9.8536e-02, -4.6085e-02,  1.4373e-01, -3.6092e-02, -2.7668e-01,
          1.6622e-01, -3.6560e-02,  2.6156e-02, -1.3146e-01,  1.2968e-01,
         -9.0749e-02, -6.9367e-02,  9.7177e-02, -4.7472e-02, -4.3903e-02,
         -1.4468e-01,  5.9552e-02,  3.0910e-02, -1.6373e-02,  3.2107e-02,
          4.4506e-02, -6.1001e-02, -6.8160e-04, -1.6244e-01, -5.2226e-02,
         -5.5585e-02, -5.1076e-02, -4.7004e-02,  2.3687e-01,  1.0325e-01,
          2.5275e-02,  1.7769e-02,  6.5248e-02, -5.7165e-02,  7.6632e-02,
          9.7758e-02, -7.6330e-02, -1.1613e-01,  1.5641e-01, -1.7924e-01,
         -3.6398e-02,  1.2080e-01,  6.0690e-02,  1.0543e-01, -2.2108e-03,
         -1.7760e-02, -1.3305e-01,  9.0361e-02, -1.0986e-01, -1.8078e-01,
         -1.1734e-01,  4.0929e-02, -1.4823e-01, -1.1167e-01, -1.3125e-01,
         -1.0211e-02, -1.5435e-01, -1.6257e-01, -3.2368e-02,  1.0663e-01,
          6.0408e-02,  7.8135e-02, -1.4825e-02, -1.4553e-01, -3.6322e-02,
         -1.2706e-01, -2.4232e-02, -1.7430e-01, -2.2189e-01,  1.1294e-01,
         -3.2351e-02,  1.1006e-01, -4.1300e-02,  1.5935e-01, -9.5063e-02,
          2.1252e-02,  2.9520e-02,  1.4116e-02, -1.0387e-01,  1.8615e-02,
         -7.9189e-02,  9.2415e-02, -1.3530e-01, -3.3983e-02,  1.9318e-01,
          1.6108e-01, -8.6596e-02,  7.6949e-02,  1.0259e-01, -7.2222e-02,
          5.3684e-02,  1.9849e-01,  1.0413e-01,  1.7264e-01,  7.2889e-02,
         -1.0847e-01,  7.3982e-02,  2.5937e-01,  1.8954e-01,  5.4603e-02,
          1.4113e-01, -7.6364e-03,  2.0701e-01,  1.6226e-01,  3.2770e-02,
         -1.3473e-01, -6.3492e-02,  7.6089e-02, -1.4355e-01,  1.4213e-01,
          1.4943e-02, -1.3370e-01,  5.3635e-03,  5.6507e-02,  5.6479e-02,
          7.2578e-02, -1.0760e-02, -1.4287e-01,  1.1125e-01,  3.6179e-02,
         -7.4857e-02,  1.4842e-01, -1.0252e-03,  1.8442e-01,  3.5145e-02,
          1.1897e-01,  1.2838e-01,  7.2968e-02,  5.2220e-03,  3.8547e-02,
          4.2794e-02, -4.0110e-02, -2.5766e-02, -8.2365e-02, -2.7382e-02,
          2.0174e-02, -1.4718e-02, -1.0327e-02,  3.3078e-02, -6.6313e-02,
          7.1547e-02,  1.4610e-01, -1.2419e-01, -1.1303e-02,  1.5027e-03,
          1.2389e-01, -5.0993e-03,  5.1281e-02,  2.1027e-01,  1.2116e-01,
         -1.4795e-01, -1.2713e-01,  1.2907e-01, -1.3849e-01,  1.4187e-01,
          1.4028e-01, -6.6228e-02, -2.0660e-02,  5.0574e-02,  2.0140e-01,
         -5.7110e-02,  1.5259e-01, -8.7248e-02,  2.3356e-02,  1.4025e-01,
          1.7228e-01,  8.7697e-03, -6.4691e-02, -3.6287e-02,  1.2926e-01},
        '{ 9.2836e-03,  1.2511e-01,  2.5538e-02,  1.9982e-01,  2.0082e-01,
          9.8671e-02,  1.8064e-02,  9.7865e-02,  7.6781e-02,  2.8093e-02,
          1.6351e-01,  1.4728e-01, -5.5845e-02, -1.4239e-01, -7.1669e-02,
          4.7575e-02, -1.4637e-02, -9.2207e-02, -4.2426e-02, -2.6675e-02,
         -1.6906e-01, -1.9708e-01, -2.6195e-02, -1.3577e-01, -4.3833e-03,
         -5.3925e-02, -1.6585e-02,  1.1266e-01, -1.0899e-01, -1.2113e-01,
         -8.5769e-02,  1.7233e-02,  1.2289e-01,  4.1140e-02, -1.9208e-01,
         -2.5054e-02, -7.4829e-02, -6.8061e-02, -8.3128e-02,  1.6932e-02,
         -1.5640e-01, -6.8852e-02,  8.3898e-02,  1.0858e-01,  1.2128e-01,
         -1.1240e-01,  1.0934e-01,  1.0056e-01,  8.8399e-02, -6.7588e-02,
         -9.2670e-02, -4.1102e-02,  4.4324e-02, -6.3208e-02, -3.6932e-02,
         -3.2465e-02,  2.1100e-02, -4.1247e-02,  8.0908e-02,  5.3465e-02,
          2.6919e-02,  4.3784e-02,  7.3533e-02,  1.3840e-01, -1.6286e-01,
         -1.6845e-02, -8.9477e-02, -9.1015e-02, -7.9907e-02, -1.7978e-01,
          8.1025e-02, -4.3614e-02,  4.7665e-02, -1.2605e-01,  2.0693e-01,
         -2.5693e-02, -4.1251e-02, -9.0130e-02, -8.3008e-02, -9.5184e-02,
          8.6560e-02,  6.8631e-02, -6.3131e-02,  4.9585e-02,  7.7017e-02,
         -4.7003e-02, -3.1285e-03, -1.2893e-01,  1.4498e-01,  1.5977e-01,
         -2.5787e-02, -2.1659e-02, -5.3832e-02, -3.1600e-04, -1.3042e-01,
          4.9067e-02, -1.6815e-02, -2.1038e-02,  3.2612e-02, -6.9364e-02,
          8.4227e-02,  9.2091e-02, -9.3478e-02, -4.6080e-02,  2.6522e-02,
          6.0443e-02,  4.3493e-02,  1.0109e-01, -5.6405e-02, -3.6400e-02,
         -8.3228e-02, -4.0274e-02,  9.9817e-02,  5.5001e-02,  1.5022e-01,
          1.7604e-01,  8.2980e-02,  1.3987e-01, -6.7163e-02, -9.2292e-02,
         -5.7605e-02,  1.1085e-01, -2.6489e-02,  7.4942e-02,  9.5194e-02,
         -3.2507e-02, -1.4501e-01,  2.1842e-02,  3.1553e-02, -1.6236e-01,
          2.2364e-02,  1.3434e-01, -5.2761e-02,  1.4182e-01,  4.6817e-02,
          1.0153e-01,  2.3258e-01,  1.2004e-01,  4.2785e-02,  1.1503e-01,
          2.4750e-02,  1.8306e-01, -6.6481e-02,  1.4626e-01,  7.4122e-03,
         -9.1575e-02,  6.3837e-02, -1.2326e-01, -7.6934e-02,  6.6768e-02,
         -4.8093e-02,  1.1994e-01,  1.1097e-01, -2.4246e-02,  2.9790e-02,
          1.2896e-01,  1.7288e-01, -1.8500e-02,  4.5597e-02,  7.1458e-02,
         -4.3240e-02,  7.1177e-03, -2.3773e-02,  1.5928e-01,  4.3187e-02,
          1.9769e-01,  1.6770e-01, -9.9574e-02,  2.0521e-01, -1.1311e-01,
         -1.0999e-01,  8.2672e-02, -1.5755e-01,  1.4463e-02,  7.7364e-02,
         -3.7508e-02,  1.8396e-01, -5.4220e-02,  5.1369e-02, -7.6391e-02,
          6.3252e-02, -6.7504e-02,  1.0171e-01, -3.0447e-02,  1.4196e-01,
          1.0277e-02,  3.9274e-02, -1.5763e-01,  1.0597e-01,  6.1923e-02,
          7.8182e-02,  6.0996e-02,  3.7719e-02,  3.1683e-02, -4.0040e-03,
         -1.1624e-01, -1.3243e-01, -1.8663e-01,  1.2244e-01,  3.7112e-02},
        '{-6.7890e-02,  7.7457e-02, -1.2484e-01,  3.8926e-02,  8.2606e-02,
         -4.7374e-02,  1.9022e-01, -1.7427e-02,  1.3374e-02,  6.8615e-02,
          1.3001e-01,  2.6470e-02, -4.8215e-02,  8.7318e-02,  9.4874e-02,
          1.1573e-01,  1.3631e-01,  1.1346e-02,  1.1858e-01,  1.2327e-01,
          8.4363e-02, -1.2269e-02,  2.3589e-01,  1.2263e-01, -3.2371e-02,
         -1.3058e-02,  4.1748e-02, -1.4984e-01,  5.0036e-02,  2.0204e-01,
          9.6120e-02, -8.0204e-02,  5.9657e-02,  1.6828e-02,  3.2572e-01,
         -1.4583e-01, -2.3988e-03,  1.6892e-01,  2.2461e-01, -9.0411e-02,
         -5.2206e-04,  7.8789e-02,  3.8625e-02,  1.5883e-02, -2.8518e-01,
          1.3084e-01, -6.6931e-02, -8.5135e-02, -1.6450e-02, -2.3674e-02,
          6.9805e-02, -2.3914e-02,  1.1851e-01, -2.6893e-02, -6.0468e-02,
         -7.0464e-02, -5.2427e-02, -2.9290e-03, -1.0839e-01, -1.2476e-01,
          4.5618e-02, -1.0652e-01, -1.4433e-01, -6.9444e-02,  4.8408e-02,
         -6.4558e-02, -7.6682e-02, -9.6562e-02,  6.0777e-02, -2.6116e-02,
          8.2796e-02,  3.3307e-02, -4.0013e-02, -9.0490e-02, -1.3762e-01,
          6.9437e-02, -6.1037e-02,  5.0923e-02, -4.2327e-03,  1.8327e-03,
         -1.1279e-02,  1.8742e-02,  9.5368e-02,  1.1349e-02, -2.1499e-02,
         -7.6118e-02,  6.4428e-02,  2.7666e-02, -1.4876e-01, -2.0109e-01,
         -1.4146e-01,  3.6629e-02,  1.7513e-02,  1.3866e-01,  5.8162e-02,
         -5.9659e-02,  1.2414e-01, -2.7376e-02,  1.5708e-01,  9.1720e-02,
          3.1057e-02,  4.1256e-02, -5.6939e-02, -4.5589e-04, -6.0988e-02,
          1.3947e-01, -1.0655e-01, -7.1992e-02,  1.1268e-01, -6.8824e-02,
          1.4314e-01,  1.9267e-01, -9.7384e-02,  7.4683e-02, -1.6989e-02,
          2.8504e-03, -1.1668e-01, -7.8287e-02, -1.8943e-01,  1.1283e-01,
          5.0424e-02,  6.1905e-02, -3.6303e-02,  1.3435e-02,  6.9368e-02,
          6.2100e-02,  1.3275e-01, -8.5982e-02,  1.1493e-01, -3.8358e-02,
          9.7889e-02, -1.5667e-01, -9.7336e-02,  1.3803e-01,  1.3665e-01,
         -6.2697e-02, -6.3050e-02,  1.5666e-01,  7.6990e-03,  6.1561e-02,
         -1.2506e-02,  1.8368e-01, -1.7279e-04, -8.5560e-02, -7.6163e-02,
          7.3676e-02, -1.1025e-01, -5.3044e-02, -4.0851e-02, -3.2267e-02,
          1.0140e-01, -1.4331e-01, -2.5604e-02, -1.6900e-02,  6.8340e-02,
         -8.1439e-02, -1.3835e-02,  6.6936e-02,  3.5801e-02, -1.2635e-02,
         -4.7174e-02,  1.3451e-01,  1.5307e-01, -1.3347e-01,  6.6362e-02,
          4.2202e-02, -2.4576e-02, -8.8809e-02, -1.1370e-01, -4.4998e-02,
          1.1812e-01,  4.9017e-02,  2.4411e-02,  1.9459e-02, -7.3385e-03,
          4.1527e-02, -1.5402e-03, -3.8684e-02, -3.5074e-02,  7.5426e-02,
         -8.5426e-02,  4.7021e-02,  1.8136e-01, -1.0234e-01, -1.2961e-01,
          8.0536e-02,  9.5121e-02,  1.0802e-01, -1.5641e-01, -8.3615e-02,
         -1.1431e-01,  1.0284e-02, -7.9433e-02,  2.0586e-02,  1.6003e-01,
         -1.3871e-01, -2.6163e-02,  1.0516e-01, -1.7648e-02,  9.7090e-02},
        '{-2.2672e-03, -3.3423e-02, -4.3653e-02,  9.9407e-02,  1.2771e-01,
          2.0245e-02,  1.6659e-01, -1.9360e-02,  3.0828e-02,  8.3141e-02,
          5.6950e-02, -8.3085e-02,  5.7839e-02,  1.9348e-01,  9.8011e-02,
          1.8276e-02,  3.4121e-02,  1.4085e-01,  1.3152e-02,  1.4928e-02,
         -5.5500e-02, -1.1179e-01, -1.1017e-01, -7.4154e-02, -6.8971e-02,
          1.0777e-01, -1.6346e-01,  5.5766e-02,  3.2547e-01,  3.2070e-01,
         -1.3926e-01, -9.9358e-02,  1.9140e-01,  1.7646e-01,  2.3580e-01,
         -1.0509e-01,  1.3049e-02,  1.7869e-01,  7.6908e-02,  1.8071e-01,
          8.9618e-02,  3.4721e-02,  3.4390e-02,  8.4609e-02, -8.2328e-02,
          7.9180e-02,  2.4518e-01,  3.3910e-04,  7.5581e-02, -3.5281e-02,
          8.8681e-02,  9.3602e-02, -6.1121e-02, -3.9173e-02,  6.6121e-02,
          8.3080e-02, -3.2268e-02, -2.6566e-02, -1.1792e-01,  1.5690e-02,
          1.1169e-01,  9.4267e-02,  1.3618e-01, -8.1086e-02, -5.6867e-02,
         -1.1040e-02,  5.7648e-02,  1.1528e-01,  6.3511e-03,  1.6673e-01,
          1.4509e-01,  8.2189e-03,  1.4731e-01, -7.6075e-02,  1.4074e-01,
         -2.2261e-02, -6.8702e-02, -3.4972e-02,  1.4337e-02, -2.9071e-02,
          1.4407e-01,  8.0731e-02,  1.2778e-02, -1.3077e-01, -1.6779e-01,
         -6.4666e-02,  5.6126e-03,  8.8608e-02, -1.1453e-01, -8.8019e-02,
         -3.7616e-02, -1.4773e-01,  4.6198e-02,  1.2036e-01,  4.2259e-02,
          1.0335e-01, -3.7486e-03,  7.5885e-02, -2.3366e-02,  1.2053e-01,
          3.2138e-02,  6.7797e-02, -8.7973e-02,  2.5812e-02, -1.5963e-01,
          1.6805e-01, -6.7808e-02,  1.4409e-01,  3.1346e-02, -6.4035e-02,
          1.2542e-02,  1.2663e-01, -5.5475e-02, -6.3047e-02, -4.9078e-02,
         -1.3567e-01, -8.6710e-02, -5.4160e-02,  1.2444e-01, -1.3095e-01,
         -1.1375e-01, -3.1552e-02,  9.8741e-02, -6.7384e-02,  4.6111e-02,
          1.4234e-02, -7.3448e-03, -2.0035e-01, -1.0569e-01,  8.2927e-02,
         -2.0342e-01, -1.7437e-01, -5.6359e-02,  7.5582e-03,  7.2612e-02,
         -5.6743e-02,  8.9393e-02, -6.1303e-02, -1.5553e-02,  7.7012e-02,
          1.2468e-01, -1.8850e-02, -3.5464e-02,  2.3841e-03,  8.6914e-03,
         -1.2327e-01,  9.1702e-02,  1.0933e-01,  2.2243e-02, -1.5794e-01,
         -1.5659e-01,  5.6635e-02,  3.6170e-02, -4.2754e-03, -1.3849e-01,
          8.4526e-02,  1.5352e-01,  9.5326e-02, -5.1947e-02, -1.3532e-01,
          1.0134e-01, -1.4049e-01, -4.3335e-02, -6.4470e-03,  1.0484e-01,
          4.0142e-02, -2.2931e-02, -5.7501e-02, -9.1275e-02, -1.7240e-01,
          1.2709e-01,  3.4553e-03,  1.5919e-01, -1.7643e-02, -1.0807e-01,
         -8.6392e-02, -1.4237e-01,  6.1451e-02,  6.8913e-02,  9.9652e-03,
          8.2561e-02, -6.8672e-02,  4.8015e-02,  1.6462e-01,  4.8556e-02,
         -4.5501e-02,  1.3473e-01,  1.8501e-01,  1.2954e-01,  8.9873e-02,
         -8.3227e-02, -7.2990e-03, -7.2966e-02, -6.9389e-02, -5.5480e-02,
         -8.1947e-02,  3.2488e-02,  2.0724e-01, -9.6737e-02, -5.8831e-02},
        '{ 1.5264e-01, -1.1945e-01,  6.6619e-02,  1.7272e-01,  4.3498e-02,
         -3.0897e-02, -5.9022e-02, -3.6492e-02,  2.0448e-01,  6.1340e-02,
         -1.4615e-01, -1.4876e-01,  1.2314e-01,  3.4676e-02,  1.2284e-01,
          2.6760e-02,  1.5756e-01,  5.4252e-02, -1.4906e-01,  1.0607e-01,
          2.8070e-01,  2.7656e-01, -2.5991e-02, -2.1617e-02, -1.8457e-01,
          7.2402e-02,  7.6159e-02,  1.1735e-01,  1.1299e-01,  1.9097e-01,
         -1.3999e-01, -7.1628e-02, -2.1305e-03, -3.6564e-02,  4.3492e-02,
         -9.1771e-02, -3.1796e-02,  6.4913e-02,  2.2706e-02,  8.8682e-02,
          1.4122e-01,  1.6988e-01,  6.1071e-02, -6.6193e-02, -2.2408e-01,
          2.4687e-01,  8.6321e-02, -3.6227e-02, -6.0173e-02, -1.5594e-02,
         -1.1553e-01,  1.5505e-02, -1.4450e-01, -5.7173e-02, -4.3065e-03,
          8.3147e-03,  2.8303e-02,  7.4740e-03, -9.1699e-02,  5.7240e-02,
         -1.0577e-01, -7.4157e-02,  6.9532e-02,  3.7703e-02, -4.6508e-03,
         -6.4253e-02, -3.5649e-02,  1.1197e-01,  2.1503e-01,  1.2009e-01,
          9.9401e-02, -9.4921e-02,  1.1585e-01, -9.1935e-02, -2.0448e-01,
         -7.2787e-02, -1.7810e-02, -1.5832e-01, -1.2184e-01, -4.6115e-02,
         -1.2141e-02,  4.0086e-02, -8.0835e-02, -9.6626e-03, -7.7504e-02,
         -3.6402e-02,  5.8042e-02,  1.7079e-01, -8.0644e-02, -1.8574e-01,
         -1.4962e-01, -3.9121e-02, -1.0409e-01,  1.4323e-01, -4.5539e-02,
          1.9326e-03, -1.2257e-02,  1.7309e-03,  8.6253e-02,  1.5837e-01,
         -4.0666e-03, -1.5195e-01, -6.2649e-03, -9.2149e-02,  5.2162e-02,
          1.0319e-01, -1.2683e-01,  1.4055e-01, -2.7110e-02, -5.7068e-02,
          5.5615e-02,  9.2452e-02,  1.9999e-02,  2.7547e-02, -1.3845e-01,
          4.0785e-02, -1.2476e-01, -1.0315e-01, -1.0555e-01,  5.4538e-02,
          1.3203e-02, -1.1732e-01, -7.2431e-02, -1.0838e-01, -9.1934e-02,
          7.7353e-02,  7.9444e-02, -1.4182e-01, -1.1475e-01,  9.4699e-03,
         -1.0727e-01, -1.0046e-02, -7.5019e-02,  1.2281e-01,  1.8144e-01,
          8.8624e-02,  5.2464e-02, -5.2799e-02,  2.0668e-02,  3.1308e-02,
          1.0065e-01, -3.0373e-03,  1.3324e-01,  7.3331e-02, -6.8923e-02,
          1.0899e-01, -1.5220e-01,  3.8332e-02,  1.1803e-01, -1.7239e-01,
          3.5420e-02,  1.0038e-01, -9.4678e-02,  1.4077e-01, -9.8747e-02,
          1.1976e-02,  7.7728e-02,  1.4239e-01,  2.0823e-01,  1.4510e-01,
          5.9875e-02, -9.8705e-02,  5.3888e-02, -6.3411e-02, -1.1541e-01,
         -8.5121e-02,  3.2276e-03, -1.6809e-01, -4.3624e-02, -1.3595e-01,
          4.5644e-02,  1.2442e-01, -2.5369e-02,  8.7942e-02, -1.5977e-01,
          5.0423e-02, -2.3382e-02,  9.8776e-02,  6.6025e-02, -5.9904e-02,
          6.4498e-02, -1.1699e-01,  1.8114e-01, -4.6464e-02,  1.4822e-01,
         -2.3446e-02,  3.7711e-02,  3.9521e-02,  6.6039e-02, -6.5919e-05,
         -1.4865e-01,  1.4482e-02, -5.3055e-02,  8.2758e-02,  4.3401e-02,
          1.3331e-01, -7.2787e-02,  1.5146e-02,  6.9397e-02,  4.7592e-02},
        '{ 9.2851e-02, -3.8848e-02,  1.6429e-01,  2.1646e-02,  6.8667e-02,
          2.5253e-03, -1.0427e-01, -2.9933e-02,  1.5635e-01, -1.1469e-02,
         -9.2895e-02,  1.1555e-01, -1.8572e-02, -6.6517e-02, -1.2072e-01,
         -6.9605e-02, -3.8669e-02,  1.0707e-01,  1.0810e-01, -1.3496e-01,
          1.4163e-01,  6.9256e-02, -8.0435e-02,  1.0820e-02,  3.0956e-03,
         -7.7636e-02, -4.3672e-02,  1.1595e-02,  1.4696e-01, -1.0693e-01,
         -1.5909e-01, -1.0348e-01,  9.2986e-02, -1.1201e-02,  1.5613e-01,
          3.4307e-02, -5.2498e-02,  1.8319e-01,  1.8839e-01,  1.8050e-01,
          1.8151e-01,  7.5935e-02,  6.0553e-03,  1.4735e-01, -5.6502e-02,
         -1.2954e-02,  1.6885e-01,  1.6707e-01, -1.3184e-01, -7.2609e-02,
         -2.9118e-02, -1.1234e-01, -1.2111e-01,  6.4967e-02, -9.6592e-02,
          4.2047e-02,  3.5774e-02,  2.4469e-01,  6.2075e-02,  5.6898e-02,
          3.4100e-02, -6.1601e-02, -3.2739e-02,  1.5057e-01,  8.4512e-05,
          4.8304e-02,  2.3358e-02,  1.4344e-01,  3.8883e-02, -8.0027e-02,
         -5.2564e-02,  6.4284e-02,  2.7706e-02, -9.1229e-03, -9.4277e-02,
         -1.9649e-02,  3.6244e-03, -3.5461e-02, -1.3483e-01,  4.2455e-02,
          4.7670e-02,  8.7539e-02,  3.4219e-02,  8.5216e-02, -2.2766e-02,
          2.9888e-02,  6.1008e-02,  8.9197e-02, -1.7260e-03,  1.9578e-02,
         -3.4795e-02, -6.7020e-02,  1.7347e-02,  7.7571e-02,  7.3353e-02,
         -4.3768e-02, -3.4070e-02,  5.6924e-02,  5.7429e-02,  2.2110e-01,
          7.0098e-02, -1.3541e-01,  3.8654e-02, -1.2258e-01, -1.0051e-01,
          1.6086e-01,  1.7357e-01,  1.8896e-01,  1.5148e-01,  1.0011e-01,
         -9.1516e-02,  3.1850e-02,  8.2623e-02, -4.3276e-02,  1.3023e-01,
          9.1473e-02, -1.5460e-02, -9.3086e-03, -7.2561e-02, -1.2342e-01,
          1.4758e-01, -1.2929e-01,  4.7175e-02, -9.6613e-02,  6.5059e-02,
         -1.3160e-01,  2.0226e-02, -1.0754e-01, -4.9239e-02, -6.1899e-02,
         -6.3968e-02, -1.2405e-01,  5.6721e-02,  1.3759e-02,  1.9502e-01,
          2.0488e-02,  1.6132e-01, -2.2176e-02,  1.3176e-01, -5.9333e-02,
          3.3015e-02,  1.0326e-01,  4.8500e-02, -6.1059e-02, -7.1091e-02,
          7.0378e-02, -1.2344e-01,  6.0658e-02, -1.6891e-01, -4.8133e-02,
         -2.0717e-02, -8.3828e-02,  6.1768e-02, -7.2680e-02,  1.5899e-01,
          1.0463e-01,  4.5841e-02,  1.5294e-01,  6.3579e-02,  1.1422e-01,
          9.7039e-02, -6.2987e-02,  1.6645e-01,  2.8907e-02, -6.4878e-02,
         -8.3227e-02, -1.3720e-01, -1.6757e-01, -9.3901e-02, -1.8215e-01,
         -8.7386e-02, -1.3167e-01,  1.4009e-01, -1.7873e-01, -1.9778e-01,
          1.5628e-02, -8.8649e-02,  4.9308e-02,  7.8360e-02, -7.5768e-02,
          9.8256e-02,  1.5799e-01,  1.3076e-01,  1.7012e-01,  7.5606e-02,
          1.1454e-01,  7.5312e-02,  2.4795e-02,  2.8567e-02, -1.8817e-02,
          1.4837e-01, -9.2182e-02, -1.2065e-02,  2.0102e-02, -5.0561e-02,
          1.1303e-01, -5.6206e-02,  1.1439e-01,  6.0349e-02, -1.5825e-01},
        '{-4.8711e-02, -3.9617e-02, -5.2108e-02,  8.9368e-02,  1.8182e-02,
          5.2856e-02, -2.3517e-02,  6.2589e-02, -3.3449e-02,  1.0220e-01,
         -4.9476e-02,  1.6768e-01, -1.5639e-01, -1.8808e-01, -2.0476e-02,
         -1.0524e-01, -6.4245e-02,  5.6080e-02, -1.4378e-01, -4.1257e-02,
         -1.5757e-01,  5.6322e-02,  2.1636e-01, -5.9422e-02,  6.8156e-02,
          5.5457e-03,  1.8126e-02,  2.0556e-01,  2.8812e-02,  2.4357e-02,
         -4.6618e-02,  6.2167e-02,  2.4383e-02,  3.6133e-01,  1.2809e-01,
          1.4187e-01,  4.5067e-02,  2.8892e-02,  2.1621e-01, -6.0614e-02,
         -1.5432e-01, -2.2776e-01, -1.5693e-01, -2.5059e-02, -4.0854e-03,
         -5.0475e-02,  2.1254e-02,  4.1787e-02, -5.3451e-02,  1.3221e-01,
         -4.5494e-02, -1.0414e-01,  3.9061e-02, -1.2166e-01, -9.7913e-02,
          5.1395e-02, -2.4533e-02, -1.1080e-01, -2.6244e-02,  4.1765e-02,
          2.0415e-04,  1.1709e-01, -2.5907e-03,  4.1377e-02,  2.6352e-01,
          3.7225e-03,  1.5276e-02, -6.6709e-02, -1.0700e-01,  1.0638e-01,
          9.2904e-02,  1.9356e-01, -1.0796e-01,  4.0940e-02,  3.5793e-02,
          8.0566e-02,  2.9270e-02, -1.1468e-01, -9.1734e-02, -1.5310e-01,
         -2.7561e-02,  2.6317e-02, -7.8470e-02, -1.0214e-01, -1.8540e-01,
         -6.3169e-02,  1.1604e-02,  4.4341e-02, -2.7405e-02, -4.1137e-02,
         -7.9094e-02,  1.6988e-01, -3.5252e-02, -4.5842e-02, -4.8866e-02,
         -1.1857e-01,  3.3049e-03,  1.0413e-01, -2.9202e-02, -1.1559e-01,
         -7.3859e-02,  3.9704e-03,  6.0421e-02, -7.2697e-02, -1.4872e-01,
         -5.6732e-03,  1.0679e-01,  1.8371e-01, -1.3171e-01, -4.7698e-02,
          1.6351e-01,  4.3335e-02,  3.4760e-02,  2.5147e-02,  1.3075e-01,
          6.4863e-02, -3.1633e-02,  7.1042e-03,  9.9824e-03, -1.0132e-02,
          9.0447e-02,  1.2633e-01, -1.0479e-01,  9.0673e-04, -9.1663e-04,
          1.0758e-01,  4.5046e-02,  1.0751e-01,  2.1277e-03,  2.6090e-02,
          3.1310e-02,  3.7230e-02,  1.6982e-01,  1.7190e-01,  3.2848e-02,
          2.1917e-02, -4.4187e-02, -5.3561e-02, -2.7209e-02,  1.0589e-02,
          7.5873e-02, -7.3582e-02,  6.7579e-02,  3.9425e-02,  7.2385e-02,
          5.3654e-02,  1.2194e-01, -2.1178e-02,  1.0476e-02, -3.0078e-02,
          2.6726e-02, -1.2273e-01,  1.1933e-02, -5.9565e-02, -5.8802e-02,
         -2.7833e-02,  6.7457e-02,  8.7465e-02, -4.6501e-02, -1.3739e-01,
          4.0943e-02,  1.6784e-02,  1.9134e-02, -1.3654e-01,  1.2387e-01,
         -3.2635e-02,  1.2301e-01,  5.5335e-02, -8.2881e-02, -6.0974e-02,
          8.1520e-02,  1.3265e-01,  1.7735e-01,  9.3446e-02,  1.5966e-01,
          5.7637e-02,  8.0196e-02,  5.1372e-02,  1.2675e-01, -2.4669e-02,
          1.3856e-02, -5.6267e-02,  4.6957e-02,  1.5707e-01,  8.3641e-02,
          9.7651e-02,  1.4344e-01,  5.9845e-02, -1.7312e-01, -4.1709e-02,
         -1.1820e-01,  1.4249e-01,  3.3810e-03, -4.9857e-02,  1.5969e-01,
          2.4096e-02, -1.3989e-02, -1.8426e-02,  4.0441e-02, -2.9060e-03},
        '{-1.5323e-01,  2.1578e-03, -2.1047e-01, -2.0342e-01, -8.3608e-02,
         -8.0719e-02,  2.8237e-02, -1.3847e-01,  6.5174e-02,  1.4659e-01,
          8.5064e-02,  3.3119e-02, -9.2268e-02,  6.8042e-02,  2.6157e-02,
         -1.1982e-01,  7.8444e-02,  1.8463e-02, -5.9259e-02,  3.9230e-02,
         -1.9507e-01, -9.5915e-03,  1.6950e-02,  9.8735e-04, -1.0716e-01,
         -1.1300e-01, -2.5833e-01, -1.7655e-01,  4.4993e-02,  1.3648e-01,
         -8.9962e-02, -2.9876e-01, -2.4406e-01,  2.3991e-02,  1.4900e-01,
         -3.0334e-01, -1.4702e-01, -1.0530e-01,  6.6676e-02, -4.8191e-02,
         -1.1665e-01,  5.1315e-02, -4.1862e-02, -8.6487e-02, -1.2601e-01,
         -2.0528e-02,  1.5492e-01,  4.3555e-02,  1.7711e-01,  1.2448e-01,
         -5.8039e-02, -7.5817e-02,  1.2181e-01,  1.2820e-01, -9.0946e-02,
          1.2752e-01,  1.5971e-01,  4.3568e-03, -4.6884e-02, -7.3242e-02,
         -6.6950e-02,  7.2344e-03, -2.7151e-01,  1.5191e-01,  1.3067e-01,
          1.3206e-01,  1.7636e-01, -6.6912e-02,  1.8822e-01,  1.4026e-01,
         -2.5059e-02,  9.4807e-02,  3.7390e-02,  1.0637e-01, -3.0265e-02,
          1.8451e-01, -4.7069e-02,  1.1817e-01,  6.5914e-02,  1.3732e-01,
          6.7589e-02,  3.7975e-02, -4.5210e-02, -4.3263e-03,  1.0376e-01,
         -8.8973e-02,  1.2623e-01, -5.9977e-02,  1.2494e-01, -1.1881e-01,
         -1.2147e-01, -3.0573e-02,  5.1751e-04,  3.5456e-02,  2.7197e-02,
         -1.1135e-01,  1.2005e-01,  7.1758e-03, -8.5239e-02, -3.6079e-02,
          3.0000e-02,  2.4787e-02,  4.2331e-03,  7.1015e-02, -1.5244e-01,
         -5.5984e-03,  5.8370e-02, -9.8851e-02,  4.4796e-02, -8.7290e-02,
          1.0621e-01,  1.8077e-01,  4.9137e-02, -1.7077e-01,  8.6604e-04,
         -6.7615e-03,  8.6447e-02,  9.9657e-02, -4.8191e-02,  5.8218e-02,
          1.1254e-01, -3.6389e-02,  5.4432e-02,  8.9833e-02, -1.3189e-01,
          2.5226e-02, -2.8372e-02, -7.1881e-02,  4.9896e-02,  1.5214e-01,
         -1.7688e-01, -1.3277e-01, -2.7622e-01, -6.9560e-02, -3.9346e-02,
         -1.2169e-01,  3.9703e-02,  6.2633e-02,  3.4873e-02,  1.4161e-01,
         -6.9306e-02, -7.1385e-02, -1.7046e-01, -4.0078e-02,  1.8601e-01,
         -1.0767e-01,  1.0539e-01,  1.1618e-01,  1.2402e-01,  1.0796e-01,
         -3.4730e-03,  3.6150e-02, -4.7599e-03, -5.2323e-02,  5.4798e-02,
          2.2431e-02,  7.2869e-02,  4.0630e-02, -1.6549e-01,  4.8290e-02,
          1.3472e-01, -4.3582e-02,  7.0086e-02, -1.5078e-01,  1.4695e-01,
          9.2041e-02,  1.2336e-01, -1.2657e-01,  1.5342e-01, -4.1195e-02,
         -4.5430e-02, -8.5229e-02,  7.8374e-02,  2.4004e-02, -6.2374e-02,
         -8.8322e-02,  1.5005e-01, -1.1545e-02, -1.3547e-01,  1.2871e-01,
         -5.0904e-02, -9.2232e-02,  8.6870e-02, -7.1634e-02, -7.2417e-02,
          1.6245e-02,  1.6384e-01, -1.0916e-01,  2.2789e-02, -3.9377e-02,
         -2.3854e-02,  3.7046e-02, -1.1928e-01,  1.1054e-01,  3.8907e-02,
         -9.6986e-02, -6.8252e-02,  1.6456e-01, -3.6891e-02, -9.3645e-04},
        '{-2.3386e-02,  1.5492e-01,  4.7266e-03,  1.4478e-01,  1.4261e-01,
          5.0308e-02,  5.0124e-02,  3.0414e-03, -1.0647e-01,  6.9524e-02,
          7.0608e-02,  1.5273e-01,  9.0900e-02,  7.9274e-02,  5.8041e-02,
          2.9503e-02,  1.5238e-01, -1.1175e-01,  1.2441e-01,  5.5250e-02,
          2.2859e-01,  2.5998e-02, -1.3557e-01, -4.0565e-02, -4.7487e-02,
          9.7867e-02, -2.8417e-03,  1.3295e-02,  2.3940e-01,  2.1491e-01,
         -3.9331e-02,  1.9639e-01,  2.1376e-01, -1.2682e-01, -1.6229e-03,
         -3.6101e-02,  8.2329e-02,  1.3205e-02, -5.6862e-02,  5.8501e-02,
         -1.6458e-02,  2.2130e-01,  2.0495e-01,  1.7146e-01,  1.7112e-01,
          2.7019e-01,  3.6965e-02,  9.0352e-02,  2.1103e-02,  6.2312e-02,
         -7.9816e-02,  1.1200e-01, -4.4183e-02,  5.9913e-02,  4.7318e-02,
         -3.8583e-02, -5.2685e-02,  9.6945e-02,  9.2863e-02, -1.7926e-01,
         -1.0402e-01, -1.2073e-01,  8.0138e-02,  1.6907e-01, -2.0295e-02,
          5.5241e-02,  1.1489e-02,  5.9995e-02,  6.6558e-02,  1.0169e-01,
         -2.9874e-02,  5.0417e-02,  8.8101e-02,  1.0724e-01,  4.4543e-02,
         -7.5560e-02,  8.4663e-02, -1.4166e-01,  1.5449e-01,  9.5164e-03,
          2.7714e-03,  3.7202e-02, -9.5967e-02,  3.7978e-02,  1.0277e-02,
          3.3274e-02,  4.4823e-02,  1.0492e-01,  1.1533e-01, -1.5526e-01,
          1.1030e-01, -1.4359e-01, -2.9661e-02, -4.6736e-02, -1.4921e-01,
         -5.1035e-02,  7.3009e-02,  1.8018e-02, -5.1169e-02,  7.0783e-02,
          6.7230e-02,  1.5891e-01, -1.0563e-01, -1.5127e-01, -1.0156e-01,
         -5.8956e-02,  1.7373e-03, -1.4237e-02,  1.6778e-02,  1.2685e-01,
          9.3838e-02,  5.6815e-02, -1.0036e-01,  1.0041e-01,  1.7828e-01,
         -1.3865e-01, -8.4915e-02,  7.1070e-02,  2.0327e-01,  1.2529e-01,
         -1.3777e-01, -1.0311e-01, -5.3374e-02,  1.0326e-02,  3.5734e-02,
          1.0978e-01, -3.8273e-02, -1.1390e-01, -5.0870e-02,  2.6780e-02,
          1.5614e-01,  1.8930e-01, -9.5059e-03, -6.7595e-02, -1.1283e-01,
         -8.8232e-02,  1.9677e-01,  3.4816e-03, -4.3968e-02, -1.5951e-01,
          2.1915e-01,  6.0690e-02,  5.6231e-02, -4.6659e-02,  4.3156e-02,
         -7.9708e-02,  7.8302e-02, -2.5647e-02,  1.6344e-01,  3.6809e-03,
          6.6795e-02,  6.1314e-02,  8.5299e-02, -9.5702e-02,  5.7765e-02,
          1.1907e-01,  1.1465e-01, -1.1676e-01,  3.0539e-02, -4.3562e-02,
         -4.8991e-02,  1.0286e-01, -3.3187e-02, -4.7249e-02,  1.0648e-01,
          1.0705e-01, -5.3783e-02,  7.2838e-02, -2.1026e-02, -8.0542e-02,
         -1.4265e-01,  2.1916e-02, -2.6879e-02, -1.3621e-02, -2.9495e-02,
          4.5685e-02,  1.1605e-01, -3.9700e-02, -1.8239e-02,  9.8935e-02,
          1.2655e-01,  8.7928e-02,  1.5452e-01,  1.5134e-01, -1.0219e-01,
          1.2402e-03,  2.7403e-04, -2.3933e-02,  1.9794e-01,  8.0055e-02,
         -1.0907e-01, -1.0199e-01,  1.5188e-01,  8.5877e-02,  1.4132e-01,
         -7.9568e-02, -4.4812e-02, -1.2904e-01,  5.0714e-02, -1.1161e-01},
        '{ 8.1783e-02,  1.7605e-01, -9.9268e-02,  9.9717e-02,  6.1771e-02,
          4.4889e-02,  1.0794e-01,  5.5660e-02,  3.7410e-02, -9.4196e-02,
          2.3905e-01, -1.4259e-01, -1.9499e-01, -4.2764e-02,  5.1268e-02,
          8.6686e-04,  5.0315e-02,  1.1488e-01, -9.7347e-02, -4.1205e-03,
         -4.2159e-02,  2.9365e-02, -1.3677e-01,  1.7656e-01,  3.1287e-02,
          7.7060e-02,  1.8760e-01,  6.9079e-02, -1.2298e-01, -8.6444e-02,
          2.4257e-01,  3.4671e-01,  5.3218e-02, -2.2980e-01, -3.3514e-01,
          1.9099e-01,  2.9162e-02,  1.4726e-01,  6.1153e-02, -2.3319e-01,
          8.5745e-02, -9.0962e-02, -1.9260e-01,  1.5477e-01,  1.4287e-01,
         -2.0035e-01, -1.8083e-01, -7.2894e-02, -7.1473e-02,  1.7848e-01,
          2.9335e-02,  1.0613e-01,  2.3023e-01,  1.3855e-01, -4.9873e-02,
          4.3604e-02, -8.3842e-02,  2.1148e-02,  8.6838e-02, -1.0219e-01,
         -9.4246e-02, -1.3168e-01, -4.2577e-02,  3.4261e-02, -1.0061e-01,
          1.1266e-01, -2.4737e-02, -1.5793e-02, -9.0431e-02, -5.0424e-02,
         -5.2721e-02, -8.7929e-02,  4.5731e-02,  7.2090e-02,  9.2632e-02,
         -1.0222e-01, -9.7685e-02, -5.3884e-02,  3.4029e-02, -1.0321e-01,
         -9.3318e-02, -9.2113e-02,  8.5823e-02,  5.5112e-02,  1.3298e-01,
          7.9164e-02, -1.5352e-01,  2.8814e-02,  1.7242e-01,  1.5570e-01,
          3.5058e-03, -1.3817e-02,  1.4097e-01,  7.1238e-02, -2.5386e-02,
          4.9509e-02,  1.0176e-01, -2.9514e-02, -6.8931e-03, -1.2440e-01,
          4.1983e-02,  4.7886e-02,  6.2872e-02, -4.8818e-02, -8.1344e-02,
          2.7909e-02, -5.8842e-02,  1.2697e-02,  1.8827e-01,  1.5776e-01,
         -2.0271e-03,  5.1857e-03,  1.5076e-01,  4.1575e-02, -4.3748e-03,
         -8.9358e-02,  1.1970e-02,  1.6517e-01,  9.2225e-02, -1.2417e-01,
          3.1538e-02, -1.5278e-02, -5.4879e-03,  7.1903e-02,  3.6024e-02,
          6.1168e-02,  1.1281e-01,  1.1445e-01, -1.3894e-01, -1.5311e-01,
         -4.4037e-03,  1.9318e-01,  1.9266e-01,  1.8311e-02, -1.5118e-02,
          3.5224e-02, -1.8659e-01, -2.9520e-02, -2.6354e-02, -4.9624e-02,
         -4.6123e-02, -1.6386e-01, -1.5217e-01,  9.3651e-02, -1.9567e-02,
          5.3163e-02, -5.9372e-02,  1.1903e-01, -7.6384e-02,  7.9439e-03,
         -1.9544e-02,  5.4355e-03, -8.9963e-02, -1.4896e-02, -8.0584e-02,
         -3.7735e-02, -5.9218e-02, -4.7761e-02,  1.0320e-01,  9.3315e-02,
          7.8870e-02, -1.0450e-01,  1.1508e-01, -5.9619e-02, -1.0740e-01,
          1.0873e-01,  9.2599e-02,  1.8768e-01, -1.2580e-02,  6.5927e-02,
          6.8577e-02,  1.4507e-02, -8.0193e-02,  9.7465e-02,  1.2965e-01,
          1.0609e-01,  8.2608e-02,  1.2847e-02,  1.4251e-01,  1.0814e-01,
          8.5640e-02, -1.0767e-01, -7.6305e-02,  1.4991e-01,  3.9827e-02,
          1.5052e-01, -1.6656e-01,  1.0362e-01,  1.1239e-01, -9.4183e-02,
         -3.7158e-02,  8.9220e-02, -1.5112e-02, -2.2649e-02,  3.4151e-02,
          1.2991e-01, -2.1183e-02,  1.3982e-01,  9.0480e-03,  1.0478e-01},
        '{ 1.0144e-03, -1.6066e-03, -1.9751e-03, -2.5028e-02, -1.0927e-02,
          1.0535e-02,  4.6357e-03,  1.1900e-02,  5.2551e-02,  3.4854e-02,
         -7.9403e-03, -2.9022e-03, -1.1302e-02, -2.7979e-03,  4.4514e-02,
         -4.1534e-02, -3.2884e-02, -3.4960e-02,  1.9730e-03,  7.8777e-03,
         -6.1977e-03, -1.7265e-02,  2.9463e-02, -4.0506e-03,  2.5988e-03,
          4.1986e-03,  4.4717e-03,  4.8098e-03,  8.2723e-04,  1.8530e-03,
         -3.8275e-03, -3.3832e-03, -5.4019e-03, -4.1413e-03,  1.0512e-03,
          4.4523e-03,  4.9576e-03, -5.1293e-02,  5.0960e-02,  4.7894e-02,
         -8.4139e-04,  4.0373e-03,  2.6090e-03,  1.4527e-02, -2.6105e-03,
         -1.0357e-03, -2.5740e-02,  2.7072e-02,  7.7224e-03,  3.2022e-03,
         -4.8995e-03, -1.0287e-03, -1.1146e-02,  2.2160e-03, -3.6998e-03,
          3.4530e-03, -3.8926e-02, -2.7180e-02, -6.1698e-03, -1.2801e-03,
          3.6292e-03, -3.8612e-03,  1.2023e-02,  4.5495e-02,  2.6901e-02,
          2.8428e-02, -1.2596e-02, -1.4508e-03, -1.0719e-02,  4.0130e-04,
         -9.3959e-03, -7.0890e-03, -6.2635e-03,  3.1191e-03,  5.0960e-03,
         -1.6313e-03, -2.1599e-03, -8.1046e-03, -3.1758e-03, -4.0022e-03,
          4.4340e-03, -3.7058e-02, -4.5551e-03, -3.2157e-03, -2.6707e-03,
          7.1471e-03, -7.6687e-03,  3.2679e-05, -9.1600e-03,  1.0278e-02,
         -1.7153e-02,  6.3410e-02, -1.1597e-03,  7.6469e-03,  7.3848e-03,
         -1.2465e-02, -5.8720e-02,  1.8846e-03,  1.0075e-02,  4.8087e-03,
         -9.5035e-04, -2.3154e-03, -1.0062e-02,  3.8802e-05, -9.8186e-03,
          5.3008e-03, -3.8788e-03,  4.1049e-02, -1.1120e-02, -5.4500e-02,
          4.7448e-03, -1.0024e-02, -6.9759e-03, -1.1377e-02, -2.1980e-02,
         -1.4117e-02, -3.1500e-02, -3.5921e-02, -1.6004e-02,  2.4349e-03,
         -4.7140e-03,  2.6498e-02, -3.3351e-02, -3.0142e-03,  5.8368e-03,
         -4.9400e-03,  2.7836e-03, -1.6123e-03,  1.5729e-03, -1.3435e-03,
          3.3285e-03,  8.6806e-04, -4.7374e-03, -7.8266e-03, -3.7918e-03,
          5.4840e-03, -2.8677e-02, -4.1272e-03, -2.9725e-02,  2.3259e-02,
         -3.4554e-04, -1.1608e-02, -2.3384e-02,  9.2452e-03, -3.1653e-02,
         -2.0697e-02,  4.3450e-02, -2.0790e-02, -2.6555e-03,  4.6733e-03,
         -1.6368e-03, -1.7474e-03, -2.9133e-04, -1.9738e-02, -7.0484e-03,
          5.7307e-03,  2.0403e-02,  7.0183e-02, -2.6361e-03,  1.5765e-02,
          4.4203e-03, -2.3532e-03,  3.1548e-02,  4.9542e-02, -2.0615e-03,
          2.6376e-02, -4.7198e-03, -7.0366e-03, -3.4912e-02,  1.1823e-03,
         -5.6916e-03, -7.0962e-03,  5.1520e-02,  2.1090e-03,  5.8710e-03,
         -1.5942e-03, -6.7063e-03, -9.4746e-03, -1.2747e-02, -6.0156e-03,
          3.1171e-03, -2.2581e-02, -4.9830e-02, -5.9278e-02, -2.0304e-02,
         -2.3654e-04, -3.6620e-02, -5.3067e-03,  1.2876e-02,  2.4296e-02,
         -4.2165e-02,  2.4594e-02, -2.3195e-02, -3.5297e-03,  6.8202e-04,
         -5.0013e-02, -1.5040e-02, -5.7696e-02,  1.9462e-03,  5.1366e-03},
        '{ 4.0173e-02, -6.1176e-03,  6.3683e-02, -4.6795e-02, -8.8383e-02,
         -4.2828e-02, -1.1691e-02, -4.7410e-02, -9.6638e-03,  7.8459e-02,
          6.0082e-02,  2.2612e-02,  1.0309e-01, -3.8137e-02,  5.5177e-02,
         -3.0781e-02, -5.2317e-02,  8.3296e-02, -6.5232e-02, -1.4513e-02,
         -1.0284e-01,  1.0188e-01, -3.4166e-02,  2.6358e-04,  1.9083e-01,
         -3.5588e-02, -1.1501e-01,  4.0244e-02,  1.4683e-01,  2.5681e-02,
         -8.3270e-03, -6.0931e-02,  1.1596e-01,  5.2959e-02,  1.7730e-01,
          8.9769e-02,  2.0700e-02, -6.3963e-03, -8.2205e-02, -2.5452e-01,
         -3.0391e-02,  1.0018e-01, -2.2806e-02,  3.8307e-02,  1.1184e-02,
         -4.8164e-02, -4.2518e-02, -1.2160e-02,  1.0259e-01, -1.9789e-02,
          5.8188e-02,  6.1605e-02, -8.4933e-03, -1.9371e-02,  4.1027e-02,
         -5.8262e-02,  1.5308e-01, -8.2602e-02, -4.9808e-02,  4.3312e-02,
          4.1085e-02,  2.1002e-02, -5.0585e-02,  8.5967e-02,  1.3407e-02,
          5.4641e-02, -7.0104e-02,  5.2212e-03,  5.7705e-02,  3.0915e-02,
         -4.9077e-02,  3.5924e-02, -2.3595e-02,  1.1844e-01,  1.3595e-01,
          8.3869e-02,  8.7557e-02,  1.3846e-01,  1.7415e-02,  3.5266e-02,
          4.1685e-02,  5.9245e-02,  2.5795e-02, -6.1768e-02, -7.1888e-02,
          2.4857e-02,  2.1573e-02, -4.2006e-02,  5.6977e-02, -2.8858e-02,
          2.3368e-02, -1.0357e-01, -6.7532e-02,  1.2613e-01, -7.0550e-02,
         -1.9685e-02, -1.9940e-02,  4.8426e-02,  7.4176e-02, -3.2278e-02,
          1.8616e-01,  1.0147e-01,  2.3742e-02,  1.3772e-01,  4.5498e-02,
         -6.7785e-03,  3.9068e-02,  9.3114e-02, -1.0128e-01, -4.0742e-02,
         -4.4778e-02, -7.6297e-02, -1.7782e-01,  4.5078e-02, -1.2598e-01,
          4.4864e-02, -1.0399e-01, -6.6222e-02,  4.0421e-02,  4.4474e-02,
          1.0540e-01,  7.1949e-02, -4.7673e-02,  8.7829e-02,  7.2064e-02,
          8.6177e-02, -1.2524e-02, -7.9715e-02,  9.8063e-02,  6.0968e-02,
          1.8270e-02, -3.5873e-02,  1.0092e-01,  1.6584e-01, -4.7325e-02,
         -6.6208e-02, -2.8631e-02,  1.6985e-02,  3.9597e-03, -1.2099e-01,
          4.9516e-02, -3.7758e-02, -1.1025e-01, -1.7799e-02,  3.4596e-02,
          3.1471e-02, -2.5448e-03,  7.3961e-03,  1.3810e-02,  1.1305e-01,
          1.0094e-01,  1.1109e-01, -3.0524e-03, -1.5006e-02, -3.1990e-02,
         -2.3103e-02,  1.2527e-01, -4.2919e-02, -1.1225e-01, -1.3319e-01,
         -5.4167e-04, -1.4948e-01, -1.0448e-01, -1.5542e-02, -1.2420e-01,
         -3.6546e-02, -1.0322e-01,  2.1946e-02,  3.9948e-02,  4.2962e-02,
          7.3707e-02, -4.0887e-04,  1.1166e-02,  1.2334e-01,  9.6871e-02,
          1.6357e-01, -3.5486e-02, -4.1766e-03,  3.7447e-02,  1.0442e-01,
          3.7323e-02, -7.4483e-02, -5.0437e-02,  6.9517e-02,  1.6802e-02,
         -1.0225e-01,  1.0522e-02,  4.6611e-02, -1.6093e-01,  1.3906e-01,
         -6.6777e-02, -1.3112e-01, -7.3906e-03,  1.0524e-03,  1.5251e-01,
          5.9814e-02,  5.2083e-02,  3.0101e-02, -1.0314e-01,  1.5108e-01},
        '{ 8.4562e-02, -2.8521e-02, -9.5068e-02, -1.3427e-01, -4.6148e-02,
          1.1036e-01,  1.2849e-01,  4.3208e-02,  1.6021e-01,  8.0683e-03,
          3.3622e-02, -1.0603e-01,  1.1278e-01,  1.0045e-01,  1.4016e-01,
          4.1246e-03, -4.5239e-02,  4.5412e-02,  1.7437e-01, -2.0393e-03,
         -2.5276e-01, -2.0193e-01, -1.7561e-01,  1.2234e-01, -1.3484e-01,
          1.5596e-02, -6.5036e-02, -2.1141e-02,  1.4250e-01,  1.8933e-01,
         -3.3312e-02, -2.2617e-01, -2.3094e-01, -1.2206e-01,  1.9764e-01,
          1.1136e-01, -9.5774e-02,  7.6780e-02,  6.7294e-02, -4.6164e-02,
          2.1138e-01, -1.4040e-01, -4.4219e-02,  5.7023e-02,  1.7684e-01,
         -3.1507e-02, -1.1282e-01, -5.8173e-02, -2.9876e-02, -1.0085e-01,
         -6.4859e-02, -1.8578e-02, -1.2330e-02,  1.3382e-01,  1.4583e-01,
         -6.8129e-02,  8.9222e-02, -8.9765e-02, -1.3429e-01, -2.2466e-02,
          1.8500e-01,  1.3025e-03,  1.8515e-01, -1.0513e-02, -3.5297e-02,
          1.0421e-01,  1.1768e-01,  6.1252e-02, -6.1782e-02,  7.6928e-02,
         -5.3949e-02, -2.5227e-02,  1.5828e-01, -8.4052e-02, -1.3266e-01,
          1.5587e-01,  6.8433e-02,  9.8066e-02,  6.0919e-02,  2.7792e-01,
         -6.0676e-02, -2.2082e-02,  1.6581e-01,  1.4574e-01,  1.1500e-01,
          1.8253e-01,  1.2218e-02, -3.1618e-02, -6.9331e-04, -1.1087e-03,
          1.2497e-01,  3.4966e-02,  1.5881e-01,  2.0886e-02,  8.9956e-02,
         -4.0001e-02,  1.8656e-01,  1.1898e-01, -4.1051e-02,  1.6290e-02,
         -2.2598e-02, -1.1258e-03, -3.7745e-03, -8.5385e-02, -2.4051e-02,
          7.4466e-02,  1.2759e-01, -8.6961e-02, -1.6646e-02,  1.1967e-01,
          9.0015e-02, -1.0010e-01,  9.7892e-02,  1.1186e-01, -1.7231e-02,
         -1.0433e-01,  9.7424e-02,  8.8958e-02,  1.2975e-01,  2.8342e-02,
          7.4081e-02,  1.3044e-02, -1.0922e-01,  1.0242e-01,  8.2517e-02,
          3.1010e-02, -1.8323e-01, -7.4510e-03, -6.9781e-02,  3.7006e-02,
          3.4309e-02, -9.2221e-02, -2.3593e-01, -1.2985e-02, -5.0432e-02,
          7.6115e-02, -9.0765e-02, -7.6219e-02,  2.1863e-02,  9.8443e-02,
         -6.3958e-02,  7.9879e-02, -1.4318e-02, -1.7877e-02,  1.4320e-01,
          9.5750e-03, -2.2561e-02,  3.2556e-02, -7.2994e-02, -1.3037e-01,
         -7.5717e-02,  6.2138e-02,  5.6437e-02, -1.2771e-01,  1.1889e-01,
         -8.6181e-02,  1.3032e-01,  7.7730e-02,  4.3650e-02, -9.0587e-02,
         -3.4287e-02,  3.0577e-02,  1.2541e-01,  1.1525e-02,  6.3451e-02,
         -1.3461e-01,  1.5658e-02,  1.9071e-01,  1.7440e-01,  1.2120e-01,
         -1.4261e-01, -1.5639e-01, -6.8915e-02, -1.3351e-01,  2.8205e-02,
          5.3524e-02,  4.7059e-02, -1.1657e-01, -1.4071e-01, -3.3567e-02,
         -4.2159e-02,  4.2629e-02, -7.3590e-02, -4.1096e-02,  2.8369e-02,
         -3.7532e-02,  5.8020e-02,  8.7616e-02, -4.4700e-03, -8.1126e-02,
         -9.2363e-02,  5.7288e-02,  1.2698e-01,  2.7141e-03, -9.7256e-02,
         -1.4372e-02, -1.2543e-01,  1.5272e-01, -5.8155e-02, -2.5439e-03},
        '{ 9.0928e-02, -2.2371e-02,  5.9312e-02,  1.6059e-01, -1.2020e-01,
          5.1315e-02, -1.2849e-01,  1.6377e-01,  5.6290e-02, -9.7552e-02,
          2.1131e-02, -5.0769e-02,  2.3633e-03,  5.2246e-02,  1.0779e-01,
          1.1080e-01,  3.7185e-02,  3.4792e-02,  1.4156e-01, -9.7612e-03,
         -1.8756e-04, -1.0670e-01,  1.7795e-01,  6.5035e-02, -9.1123e-03,
         -6.5263e-02, -1.4331e-01, -1.1008e-01,  1.9000e-01,  2.9039e-01,
          6.5953e-02, -1.8759e-01, -1.4000e-01,  1.0003e-01,  1.1059e-02,
          2.0352e-01,  8.1391e-02, -1.3934e-01,  5.6779e-02,  1.6149e-01,
          1.1209e-01, -1.1321e-01,  9.5050e-02,  3.9750e-02, -3.5520e-02,
         -1.1137e-01,  1.2300e-01,  1.9718e-02, -2.0959e-01, -1.0894e-01,
          1.3350e-01,  1.1363e-01, -3.2397e-02,  1.8827e-02,  1.0331e-01,
          1.6145e-01, -8.1339e-02,  1.4861e-02, -1.8828e-01, -1.9418e-02,
          1.3566e-01,  2.0471e-01,  1.6236e-01, -2.8935e-02,  9.9365e-02,
          3.8958e-02, -1.0008e-01,  7.4618e-02, -1.4309e-02,  2.0853e-02,
          7.5008e-02, -7.6680e-03, -9.5464e-02,  1.4206e-02,  4.4821e-02,
         -5.5811e-02,  4.5172e-02,  1.2622e-01, -2.0378e-03,  2.4610e-02,
          4.8119e-02,  1.3166e-01,  6.9923e-02, -1.7058e-01,  3.4566e-03,
          1.1849e-01,  4.1240e-02, -7.7406e-02, -1.8828e-01, -1.2660e-01,
          2.9312e-02,  1.0820e-01,  1.7292e-01, -8.7114e-02,  6.5395e-02,
          3.0021e-02,  1.5033e-01, -5.4627e-02, -3.1663e-02,  5.3202e-03,
         -1.2301e-01, -8.8198e-02,  1.5805e-01, -1.0221e-01, -8.4065e-02,
          3.5173e-02, -1.0731e-03,  1.6583e-01,  3.4821e-02, -1.6007e-01,
          3.2949e-02,  1.2114e-01, -2.9002e-02,  3.9102e-02,  8.8053e-03,
          7.0791e-02,  8.7480e-02,  1.2935e-01,  7.5842e-02, -1.8227e-01,
          1.3318e-01,  7.9204e-02, -2.5463e-02,  7.1399e-02, -3.9601e-02,
          9.1465e-02, -1.1306e-01,  6.3469e-02,  1.3719e-01,  1.3190e-01,
         -8.5235e-02, -1.4083e-02, -1.1082e-01,  2.0071e-02,  1.2028e-01,
         -4.2636e-02,  3.6053e-02,  8.6083e-02, -1.1967e-02,  1.9844e-01,
         -6.2289e-02, -5.3185e-02,  1.6005e-01,  3.6144e-02, -1.5044e-01,
         -3.3697e-02,  7.3551e-02, -1.8417e-02,  4.0412e-02, -4.9905e-02,
          1.2657e-01,  5.0526e-02,  1.5135e-01,  3.7813e-03, -1.2121e-01,
          1.3489e-01, -7.1202e-03, -2.0735e-02, -3.1085e-02,  6.7677e-02,
          3.2765e-02, -3.0590e-02,  9.4207e-02, -1.3387e-02, -1.4789e-01,
         -4.1595e-02, -6.6648e-02,  1.0918e-01, -7.2851e-02,  8.4355e-02,
         -6.0555e-02, -1.0874e-01,  6.9876e-02,  3.6212e-02,  1.0490e-01,
         -9.7957e-02,  1.4632e-01,  1.2012e-01,  1.1782e-01, -6.7492e-02,
          2.3212e-03,  6.4418e-02, -1.9929e-02, -1.3551e-01, -1.0711e-01,
         -1.0805e-01, -3.1424e-02, -8.9626e-03,  1.1485e-02, -1.6945e-01,
          3.6208e-02, -6.0437e-02,  1.0244e-03,  1.3235e-01,  6.9045e-02,
          1.3762e-01,  1.3844e-01, -6.3727e-02,  1.8155e-01, -2.8499e-02},
        '{ 1.4302e-01,  1.2997e-01,  7.8552e-02, -1.3346e-01,  1.3047e-01,
          1.4942e-01,  4.8345e-02, -1.6796e-03,  1.5894e-01,  1.3809e-01,
         -1.0002e-01, -1.5906e-01, -2.7422e-02,  1.1139e-01,  1.1780e-02,
          1.5136e-01,  1.1082e-01, -1.1252e-01, -1.2369e-02,  1.5493e-01,
          3.6296e-02,  9.0264e-02,  6.5584e-02, -5.2407e-02, -5.4927e-02,
         -8.8783e-02, -4.5538e-02,  2.2268e-01,  7.6545e-02,  4.8508e-02,
         -8.0301e-03,  2.2957e-01,  8.6560e-02,  6.8345e-02,  1.5650e-01,
          3.8768e-02,  1.3920e-02, -6.8173e-02,  1.8700e-01,  1.6544e-01,
          1.0003e-01,  2.7782e-01, -8.2497e-03,  4.0187e-03, -1.0274e-01,
          2.2107e-01, -2.8293e-02,  3.6180e-02,  1.2812e-01,  1.4723e-01,
          5.4440e-02, -1.1411e-01, -1.6416e-01, -4.4229e-02,  3.5204e-02,
          1.4492e-01, -2.3015e-02, -9.5320e-02, -1.7806e-01,  9.2456e-02,
         -1.2437e-01, -1.4568e-01, -1.4495e-02,  6.3408e-02,  1.0989e-01,
         -1.7599e-02, -8.7163e-02,  1.2663e-01,  1.4973e-01, -4.1901e-02,
         -4.4010e-02,  2.4644e-03, -2.6545e-02, -1.6567e-02,  2.1414e-02,
         -3.0263e-02,  6.1362e-02, -1.7340e-01, -2.7262e-03, -9.0886e-03,
         -1.1710e-01,  2.8324e-02, -1.6950e-03, -1.5118e-01, -3.2603e-02,
         -7.1173e-02,  1.0045e-01,  1.6826e-01,  8.7849e-04, -2.3059e-01,
          3.1209e-02,  1.7804e-02,  5.3737e-02, -4.3407e-02, -2.5486e-02,
          4.7494e-02, -8.8585e-03, -7.7929e-02,  5.7444e-03, -3.3409e-02,
          1.8775e-01, -9.3223e-02, -2.6845e-02,  3.7586e-02, -1.3304e-01,
         -2.2944e-02,  1.0274e-03,  5.8076e-02,  7.2803e-02,  7.3224e-02,
         -1.0961e-01, -6.9959e-02,  4.6706e-02, -1.2701e-01,  1.1468e-01,
         -6.7582e-02, -2.3956e-02, -7.9944e-02, -3.9090e-02,  1.6523e-01,
          7.5348e-02, -1.1610e-01, -9.4318e-03,  7.5003e-02, -2.2451e-02,
          7.7420e-02,  1.7539e-01,  2.3223e-02, -4.7533e-02,  1.3341e-01,
          1.0729e-01,  7.6162e-02,  8.0600e-02,  5.8211e-02,  2.0759e-01,
          1.0941e-01, -1.2232e-01, -9.2777e-02,  7.4344e-02,  1.1700e-01,
          1.6715e-02,  1.1950e-02, -7.3795e-02, -8.1489e-02, -1.0582e-01,
          1.6247e-02,  1.3996e-02, -2.7139e-02, -4.5550e-02,  4.9148e-02,
          7.9529e-02,  1.5986e-01, -1.4189e-01, -1.4097e-01,  4.5302e-02,
          2.8549e-02,  3.1154e-02,  5.8192e-03,  1.5031e-01,  4.9812e-02,
         -1.0929e-01,  9.5181e-02, -9.4731e-03,  9.0867e-02, -4.9250e-02,
         -1.2150e-03, -1.4502e-01, -1.8428e-01, -1.0633e-01,  7.0480e-02,
         -3.6387e-02,  1.0296e-01,  4.1724e-02, -2.3914e-02, -6.5792e-04,
         -5.9509e-02,  1.3668e-01, -7.1989e-02, -1.1043e-01, -2.9255e-02,
         -3.0050e-03, -4.6073e-02, -1.9129e-02,  1.6392e-01, -6.4020e-02,
         -3.4464e-02, -7.8589e-02,  9.6945e-02, -2.2435e-03,  7.4223e-02,
          1.1378e-01, -9.9603e-02,  1.7157e-02, -2.1265e-02,  7.2528e-02,
         -9.9691e-02,  1.3513e-01,  1.6016e-01,  5.8911e-02,  5.8835e-02},
        '{ 1.0496e-01,  5.4604e-02,  3.2012e-02,  5.3087e-02,  1.4332e-01,
         -5.2157e-02,  1.2493e-01, -2.7511e-02,  1.1139e-01, -4.8930e-02,
          2.5522e-03, -4.8033e-03, -8.7595e-03, -9.7641e-02, -1.6311e-01,
          1.9349e-01,  8.3097e-02,  2.6508e-02, -1.2293e-02,  1.0176e-01,
          1.0939e-02,  1.9682e-01,  1.8116e-01,  1.4232e-01,  4.6779e-02,
          1.1808e-01,  1.6216e-01,  1.5344e-01, -2.3956e-01, -2.3936e-01,
          1.8573e-01,  1.2817e-01,  1.2878e-01, -1.9452e-01, -2.4839e-01,
          1.1238e-01,  4.8974e-02, -1.5442e-01,  2.1303e-03,  3.5552e-01,
          1.1871e-01,  4.2747e-02,  1.9099e-02, -4.7500e-02,  8.9660e-02,
          7.5970e-02,  6.4333e-02, -2.2503e-01, -1.6946e-01, -9.4945e-02,
         -1.2199e-01,  5.8591e-02,  4.0692e-02,  5.0551e-02,  3.4539e-02,
         -7.7856e-02,  1.4491e-01,  1.1389e-01, -1.6001e-02, -1.0427e-01,
          2.9658e-02,  2.0134e-01,  2.3258e-02, -8.3647e-03, -1.6698e-02,
         -5.5115e-02,  1.8574e-02,  1.5694e-01, -5.4980e-02,  1.4647e-01,
         -4.6675e-02, -1.7196e-01, -8.7504e-03,  1.4881e-02, -1.1436e-02,
         -3.2810e-02, -1.5752e-02, -5.6517e-02,  4.4234e-02, -2.1758e-01,
         -3.4768e-02,  2.5457e-02,  8.5590e-04,  6.3475e-02,  2.6588e-02,
         -4.0103e-02,  2.9328e-02, -1.6628e-02, -8.1458e-02, -1.5765e-01,
          2.6499e-02, -3.1321e-02,  5.9377e-02, -1.8129e-01,  2.2160e-02,
         -2.5669e-03,  5.8248e-02, -5.2799e-02, -1.0994e-01,  2.8424e-02,
          5.4485e-02, -3.4138e-02,  2.2993e-01,  2.1616e-01,  1.8571e-02,
         -1.3479e-01, -1.8450e-01,  2.7617e-02, -1.0670e-01,  1.3714e-01,
          7.9593e-02,  9.2399e-02, -1.1877e-02,  1.4863e-01,  1.7456e-02,
         -1.0506e-01, -3.7537e-02,  1.1594e-01,  3.5977e-02, -1.1860e-01,
          2.2069e-01,  8.8044e-02,  1.5580e-01, -1.2236e-02,  2.0217e-01,
         -6.2582e-03,  4.9913e-02,  1.5043e-01,  8.3886e-02, -1.7824e-01,
          1.9802e-01,  1.7878e-01, -2.4808e-02, -5.4382e-02, -1.1795e-01,
         -9.2378e-02,  6.6962e-02, -9.0304e-03,  1.6036e-01,  1.2536e-01,
         -1.7312e-01, -5.6613e-02,  1.3563e-01,  1.0395e-01, -1.5750e-01,
          5.0302e-03,  4.1876e-02,  3.8969e-02,  1.1273e-01,  1.8122e-01,
         -8.1877e-02,  1.2432e-02,  7.9994e-03, -5.7320e-02,  1.0099e-01,
         -8.1003e-03, -1.9338e-01, -7.3594e-02, -7.4514e-02, -4.9533e-02,
         -5.1057e-02,  1.4943e-02,  1.7992e-01,  4.7228e-02,  3.8836e-02,
         -2.6631e-02, -2.4596e-02, -1.0490e-01,  3.2882e-02,  1.1307e-01,
          6.9283e-02,  1.3221e-01,  5.5486e-02,  1.5255e-01,  2.4764e-01,
          2.5654e-02,  5.0745e-02,  7.2338e-02,  1.5104e-02,  1.9452e-01,
          2.4076e-04,  1.5417e-02, -6.9441e-02,  2.3024e-03,  1.6909e-02,
          2.4734e-02, -6.3482e-02,  1.9659e-01, -6.6564e-03,  4.7578e-02,
          3.9456e-02, -1.3643e-01, -4.2997e-03, -4.3620e-02, -1.2988e-01,
          5.1214e-02,  4.3646e-04, -5.6198e-02,  9.7516e-02,  1.2599e-01},
        '{-5.1083e-02, -1.0545e-01, -4.4256e-02,  4.9556e-02,  1.1100e-01,
          1.1813e-01,  5.0475e-02, -6.2464e-02,  6.7800e-02,  1.0997e-01,
         -8.5112e-03,  4.2022e-02,  1.5275e-01,  1.7794e-01,  5.0547e-02,
         -6.0797e-02,  1.5025e-01,  2.0212e-02, -2.5624e-02, -1.2970e-01,
         -4.6142e-03, -2.0827e-01, -6.2136e-02, -1.0627e-01, -1.1634e-01,
         -1.4685e-01, -2.1498e-01,  2.6981e-02,  1.4337e-02,  1.4639e-01,
         -2.0315e-02, -2.6680e-01, -2.2596e-01,  3.1143e-04,  2.2047e-02,
         -2.8494e-01, -2.8369e-01, -1.2780e-01, -2.7363e-01, -4.5803e-02,
          7.9063e-02, -1.0781e-01, -8.9640e-02, -9.6286e-02,  4.7055e-02,
          9.3003e-02, -1.4667e-01,  9.5725e-02, -1.4853e-01, -3.6819e-02,
          1.1515e-01,  1.3309e-01,  1.2268e-01,  1.1493e-01,  5.4787e-02,
          3.1469e-02,  1.7969e-01, -5.2843e-03,  6.7310e-02,  5.3328e-02,
         -1.2200e-02, -1.1535e-01,  8.5556e-02,  1.9525e-02, -1.2525e-01,
          1.5403e-01,  1.6768e-01,  1.0255e-01, -4.2130e-02,  4.0202e-02,
         -7.7796e-02,  1.1071e-01,  2.1619e-01, -1.7421e-02, -1.1162e-01,
          5.0626e-02,  1.1516e-01,  1.9858e-01,  2.1150e-01,  1.7478e-01,
          1.2877e-01,  9.9803e-02,  1.4062e-01,  1.7198e-01,  7.9277e-02,
          9.1898e-02,  1.2730e-02, -4.6910e-02, -2.8658e-02,  1.6110e-01,
          3.4858e-02, -1.6744e-02, -2.2631e-02, -1.6835e-02, -2.3213e-02,
          8.1573e-02, -7.9385e-03, -1.0883e-02, -1.2602e-02, -5.6908e-02,
          1.5043e-01,  1.4482e-01,  5.1057e-02,  2.1811e-02, -1.0416e-01,
          8.8495e-03,  7.9264e-02, -1.2587e-01, -6.0822e-02, -4.3916e-02,
          8.8625e-02,  1.0958e-01, -1.2113e-02,  2.0600e-01,  1.7669e-01,
          5.0532e-02,  2.9782e-02, -6.1037e-02,  1.4959e-01,  9.8325e-03,
          3.7575e-03,  9.2221e-02, -1.2198e-01,  5.4926e-02, -1.4577e-01,
          9.3513e-02, -3.0730e-02, -1.0698e-02,  1.1550e-02,  1.4045e-01,
         -1.7771e-02, -2.8202e-02, -1.2327e-01, -2.4886e-01, -9.2052e-02,
         -1.2412e-01, -4.5869e-02, -1.5278e-01,  3.8088e-02,  9.3941e-02,
          8.7861e-02, -1.0317e-02, -2.8774e-03, -5.2138e-02,  9.3603e-02,
         -1.8911e-01,  6.1663e-03, -9.7487e-02,  5.3180e-03, -1.1998e-01,
         -1.0703e-01,  1.4358e-01,  1.6195e-01,  1.1482e-01, -1.2827e-01,
         -5.8952e-02,  1.7292e-01,  1.1987e-01, -1.3595e-01,  5.8712e-02,
          1.1690e-01,  7.4811e-02,  5.2932e-02, -7.2847e-02,  1.0430e-01,
          7.5911e-03,  2.4557e-02, -1.0139e-01, -5.3066e-02,  7.4727e-02,
         -1.2640e-01,  1.6564e-02, -6.4734e-02, -8.4848e-02,  3.8672e-03,
          1.6208e-01,  1.3043e-01, -1.1544e-01,  7.3854e-02,  2.8557e-02,
         -7.7070e-02,  5.4567e-02,  1.3560e-01, -9.0176e-02,  1.3522e-01,
          8.8089e-02,  4.1239e-02, -1.5467e-02,  4.3566e-02,  1.1668e-01,
         -3.9450e-02, -6.0199e-02, -8.7576e-02,  7.2657e-02,  5.0831e-02,
          4.9734e-02, -1.6865e-01, -4.0062e-02,  1.0276e-02, -1.0093e-01},
        '{ 6.7375e-02,  1.6665e-03, -5.8992e-02,  8.5949e-03,  1.0144e-01,
         -6.0855e-02, -4.5453e-02, -1.1248e-01,  6.9222e-02, -1.8186e-01,
          1.0521e-01,  2.2566e-02,  1.1813e-01, -1.4246e-03, -2.3789e-02,
          8.9997e-02,  4.5804e-02,  7.5879e-02,  3.7572e-02,  7.3476e-02,
          7.0587e-02, -2.0465e-02,  2.1435e-01,  1.1390e-01,  4.3741e-02,
          1.1373e-01,  8.1859e-02, -1.1356e-01,  2.5103e-02,  2.4161e-01,
          1.5804e-01,  2.4040e-02,  9.0166e-02, -2.8488e-03,  8.2353e-02,
          1.7279e-01, -8.3233e-02, -2.1541e-01,  2.0804e-01,  1.4540e-01,
          6.1895e-02, -1.3631e-01, -1.5291e-01,  2.7221e-02, -4.2347e-02,
         -1.3848e-01,  4.4066e-02,  8.6161e-02,  7.2671e-02,  2.6083e-02,
          1.2713e-02,  1.2658e-01,  8.4786e-03,  1.5878e-01,  1.1796e-02,
          1.3493e-01, -3.5355e-02, -1.1592e-01, -7.5323e-02, -8.0580e-02,
          5.9868e-02, -5.0527e-02, -1.6203e-01, -1.3946e-01,  2.3464e-01,
          1.5668e-02,  9.3650e-02, -1.4779e-01, -1.8350e-01,  1.0635e-01,
         -7.6547e-02,  4.6992e-02,  8.5893e-02,  1.4246e-01,  7.5445e-02,
         -4.6454e-03,  1.2333e-01,  1.1914e-01,  2.2472e-01,  2.6391e-01,
         -3.6487e-02,  6.2249e-02,  1.7207e-01,  1.5851e-02,  1.5858e-01,
          1.1191e-01,  3.0730e-04,  1.1375e-01, -4.0470e-02, -2.4879e-02,
         -9.9593e-02, -9.3580e-04,  1.1104e-01, -5.1717e-02, -9.6428e-02,
         -8.8926e-02, -1.3957e-02, -1.2099e-01, -1.7395e-01, -5.9805e-04,
         -8.2618e-02,  1.2898e-01,  4.4358e-02,  1.8919e-01, -7.2547e-02,
          4.0944e-02, -1.4570e-01,  1.4871e-02, -7.1266e-02,  7.0952e-02,
          1.4574e-02,  1.0360e-01,  1.6867e-01,  1.0331e-01,  2.9768e-02,
         -7.6263e-02,  1.5672e-01,  1.9205e-01,  1.4162e-01,  8.7202e-02,
          7.6171e-03, -2.9322e-02,  2.1753e-01,  1.8421e-01,  2.3165e-01,
          6.7230e-02,  2.0881e-02, -6.6581e-02,  1.7502e-01,  1.6117e-01,
          1.7035e-01,  1.7450e-02, -2.3530e-03, -2.4308e-02, -3.0662e-02,
         -1.6089e-02, -3.0646e-02, -9.3378e-02, -9.8812e-02,  1.2066e-01,
          5.9272e-02,  6.0106e-02, -8.1760e-02, -7.5982e-02, -1.9333e-02,
          1.0994e-02,  1.4419e-01,  2.2501e-01, -8.0467e-03,  3.5997e-02,
          1.2217e-01,  5.0892e-02,  6.1726e-02, -1.5074e-02, -1.3184e-01,
          6.2814e-02, -7.8513e-02,  1.2466e-01, -2.0625e-01, -1.3591e-01,
          1.4371e-01,  9.8813e-02,  1.3073e-01, -1.8178e-01, -1.0334e-01,
          6.2087e-02,  3.5472e-02,  9.4820e-02, -1.1429e-01,  3.3381e-02,
          1.4063e-01,  4.5341e-02,  1.8620e-01,  7.1409e-02,  1.2852e-01,
         -7.4054e-02, -9.4124e-02,  7.7404e-02,  3.8920e-02, -1.1481e-01,
          2.9823e-02, -1.3375e-01, -7.2913e-02, -5.7881e-02, -1.0553e-01,
         -1.3503e-01,  8.1490e-02, -2.2048e-03, -5.1003e-02,  1.2826e-01,
          7.0134e-02,  2.2549e-01, -5.4065e-02, -1.3884e-01,  3.4234e-02,
         -6.5137e-02,  5.5303e-02,  4.9410e-02, -1.9205e-04,  1.6940e-01},
        '{-1.2023e-01, -1.0102e-01, -2.9454e-03,  8.0630e-02,  4.7672e-02,
          1.1171e-01, -7.2771e-02, -3.1443e-02, -3.1778e-02,  7.9516e-02,
         -5.2619e-02, -3.4514e-02,  1.3891e-01,  2.2609e-02,  2.0207e-01,
         -6.3242e-02,  2.2235e-02,  6.5258e-02, -1.2778e-01, -4.5770e-02,
          2.8044e-03,  7.9266e-02,  9.5299e-02, -1.4828e-01, -2.2553e-01,
          8.0838e-02,  6.8303e-02, -1.2228e-01, -1.8363e-01, -2.9140e-01,
         -1.4596e-01, -7.1903e-02, -2.0798e-01, -2.3495e-01, -1.7360e-01,
         -2.0080e-01, -2.7110e-01, -1.9070e-02, -8.5761e-02, -3.6392e-02,
         -4.3886e-02,  5.4903e-02, -1.3387e-01,  3.2750e-02, -4.2641e-02,
          1.3796e-01,  6.7992e-02, -7.0061e-03, -5.5612e-02, -1.8213e-01,
         -3.6354e-02,  5.5826e-03,  6.5336e-02,  7.3934e-02, -9.2573e-03,
         -1.0010e-02,  4.2866e-02, -8.8321e-02,  3.8775e-02, -9.0482e-02,
          6.1207e-03, -1.0648e-01, -2.0971e-01,  7.1439e-02, -6.4050e-02,
          6.8512e-02, -2.5393e-02, -3.9914e-03,  1.5195e-02,  6.2537e-02,
         -4.9034e-04,  3.9377e-02,  7.8901e-02,  1.9661e-02, -3.6476e-03,
          7.8279e-02, -6.5558e-02,  1.4966e-01,  1.4702e-02,  7.2780e-03,
         -5.5355e-02,  1.6618e-01,  4.2587e-02,  1.0294e-01,  8.3455e-02,
          4.3192e-02,  2.6703e-02, -7.0663e-02,  1.0659e-01,  1.2535e-01,
         -6.7902e-02,  5.0075e-03, -9.5579e-02,  1.0236e-01,  1.2720e-01,
         -1.7402e-01,  4.7748e-02,  3.3929e-02, -1.4303e-02,  1.4282e-02,
          4.6641e-02, -1.3193e-02,  3.9426e-02, -1.0088e-01, -5.9191e-03,
          1.4410e-02,  4.1897e-03, -8.3608e-03, -5.0256e-02,  3.8521e-02,
          5.3632e-03,  1.5090e-01,  8.6916e-02, -4.1402e-02, -1.3078e-02,
          1.0074e-01, -2.2571e-02, -1.7268e-01, -5.7991e-02,  6.5174e-02,
          5.8686e-02,  7.1599e-02, -1.4231e-01,  1.5101e-01,  5.3554e-02,
         -2.9875e-02, -6.4186e-02, -3.1294e-02, -1.3723e-01, -9.2577e-02,
         -1.0069e-01, -1.8572e-01, -1.7153e-01,  1.3346e-01, -1.1949e-01,
         -1.8271e-01, -2.2256e-02,  1.2603e-04, -3.6849e-02, -8.6104e-02,
          1.5053e-01,  1.8334e-01,  1.2914e-01, -8.3841e-03,  5.2312e-02,
          3.7220e-02,  1.1507e-01, -9.5528e-02,  1.5214e-02, -1.1000e-01,
          1.2935e-02,  5.9449e-02,  1.4040e-01,  3.8669e-02, -4.2333e-02,
         -4.6952e-02, -5.5624e-02, -5.3935e-02, -9.8535e-02, -4.2361e-02,
         -6.7860e-02,  4.2153e-02, -3.9721e-02,  1.3817e-01,  1.7204e-01,
         -5.8889e-02, -1.4941e-01, -1.0221e-01, -6.8476e-02,  1.7725e-01,
          9.3465e-02, -1.1299e-01,  3.9632e-02,  1.5077e-01,  5.3203e-02,
          5.8544e-03, -1.1214e-01, -2.3762e-03,  3.5738e-02, -6.0799e-02,
          6.8888e-02,  1.4851e-01,  9.5177e-02,  1.4875e-01,  2.1126e-01,
          1.6934e-01,  1.3253e-01,  3.7128e-02,  1.2414e-01,  1.6769e-01,
         -1.4475e-02,  3.3775e-02,  4.7056e-02,  1.3839e-01,  1.8206e-01,
          1.7619e-02, -7.4586e-02, -7.1510e-02,  1.1305e-01, -7.5869e-02},
        '{ 3.7442e-02,  1.2894e-01,  9.6741e-02,  1.3094e-01, -6.3900e-02,
          5.4169e-02,  5.5114e-02, -6.7688e-02,  1.9745e-01,  1.1677e-01,
         -1.0203e-01, -1.3575e-01, -2.8707e-02, -1.1234e-02,  1.0247e-01,
         -1.0389e-02,  5.1021e-03, -1.3770e-01, -4.3615e-02, -1.5622e-01,
         -1.3987e-02, -1.5582e-01, -1.4554e-01, -1.7543e-01, -1.7159e-03,
         -7.4237e-02,  2.5886e-01, -6.2707e-02,  4.5397e-02,  3.6254e-02,
         -1.0437e-01, -3.9054e-02,  2.6913e-01,  9.9177e-02, -2.0973e-01,
          8.0286e-02,  6.0353e-02,  1.7938e-01, -1.2111e-01,  6.4615e-03,
          1.6408e-02,  1.4247e-02, -4.4010e-02,  6.0291e-04,  5.1618e-02,
         -1.0569e-01, -1.3969e-02, -5.3268e-02,  2.5617e-02, -1.7435e-01,
          8.6009e-02, -1.8277e-01, -1.6454e-01, -1.8378e-01,  1.9383e-03,
          9.6355e-03, -1.1384e-01,  2.5526e-02,  2.4071e-01, -2.6359e-02,
          1.0532e-01, -8.6090e-02, -2.9541e-02, -3.7524e-03, -2.7690e-03,
          1.5801e-01, -5.9126e-02, -1.0498e-01,  6.7514e-02, -1.3192e-01,
         -1.4455e-01,  3.9101e-02,  1.6232e-01, -6.4822e-03,  1.3266e-01,
         -1.6552e-01, -7.9208e-02, -8.3436e-02, -1.4586e-01, -1.0351e-01,
         -4.6508e-02, -1.4268e-02, -1.7395e-01, -5.6622e-02, -7.9795e-02,
          1.4436e-01, -6.3646e-02, -2.7696e-02,  2.1693e-02,  1.6871e-01,
          1.2713e-01, -1.8189e-02,  6.7838e-02,  5.5270e-02, -3.2620e-02,
          7.1725e-02, -1.1553e-01, -3.5957e-02,  4.1836e-02,  2.7569e-02,
         -9.9388e-02,  9.3039e-02,  8.8480e-02,  9.2446e-02, -1.4792e-01,
          1.5985e-02, -3.9545e-02,  8.0363e-02, -5.1450e-02, -1.4408e-02,
          4.6095e-02, -1.5644e-01, -1.5228e-01,  7.0995e-02,  1.1374e-01,
         -1.4929e-01, -8.6899e-02, -9.8361e-03,  1.9393e-01,  9.5757e-02,
         -8.5274e-02, -1.2328e-01,  8.1063e-02, -8.4819e-02, -1.5411e-02,
         -1.4030e-01, -1.1796e-02, -1.1763e-01, -4.5228e-02, -5.7330e-02,
          6.5750e-02,  5.4765e-02,  2.1253e-01,  1.6905e-01, -5.7910e-02,
          6.1732e-02,  5.7242e-02,  9.1613e-02,  1.2331e-01, -8.2276e-02,
         -8.8031e-02, -7.6816e-03, -3.1498e-02,  1.1135e-01, -1.7158e-01,
          1.8042e-02, -1.6315e-01, -9.1707e-02, -1.6417e-01, -1.7466e-01,
         -1.2674e-01, -6.2687e-02, -3.5469e-02, -7.6386e-02,  1.3411e-01,
          7.0291e-03, -4.7677e-02,  4.1321e-02, -5.1387e-02,  1.3750e-01,
         -1.3542e-01, -1.6992e-01, -6.9690e-02,  1.5441e-01,  2.7887e-02,
         -7.9189e-02,  6.7847e-02,  2.0436e-01,  9.7800e-02, -1.2188e-01,
         -5.1091e-02,  5.0248e-02, -6.0865e-02,  1.3474e-02, -1.5731e-01,
         -1.4920e-01, -1.6178e-01, -4.3462e-02, -1.3866e-02,  9.8747e-02,
          3.5588e-02,  8.1442e-02,  9.7925e-04,  1.9142e-01,  1.5288e-01,
          2.9370e-02,  6.7751e-02, -3.1614e-03,  2.2881e-02, -8.7941e-02,
          8.6954e-02, -1.5875e-01, -8.6932e-02,  1.3795e-01,  4.8171e-02,
          8.0198e-03,  3.5052e-02, -3.5880e-02,  1.2071e-01, -1.7745e-01},
        '{ 8.0066e-03, -8.2132e-02,  1.8333e-02, -6.6011e-03,  5.3295e-02,
         -3.5717e-02,  1.4746e-01, -8.2507e-02,  1.3498e-01, -5.0978e-02,
          5.3016e-02,  1.0040e-04,  1.2904e-01,  1.3871e-01,  4.5071e-02,
          2.2839e-01, -1.1631e-02, -9.1912e-02,  1.1439e-01, -5.0860e-02,
          5.9796e-02,  1.4699e-01,  2.3629e-01,  1.1869e-01, -2.5084e-02,
          6.3408e-02,  1.1865e-01, -3.7102e-02, -4.8827e-02, -2.7432e-01,
         -6.4564e-02,  1.3582e-01,  1.0253e-01,  4.1524e-02, -2.7418e-01,
         -2.2322e-02,  2.1663e-03, -6.7537e-02,  7.4022e-02,  1.0763e-01,
          9.2511e-02, -8.1162e-04,  1.3102e-01, -1.8346e-02, -1.8009e-01,
         -2.8497e-02, -2.4794e-02, -2.9951e-03,  7.1233e-02, -2.3019e-02,
          4.9063e-02, -1.6404e-01, -1.3464e-01, -3.8215e-04,  1.9768e-02,
         -1.5103e-01, -1.3797e-01,  2.0463e-01,  1.6186e-01,  2.7963e-02,
          4.1492e-02, -1.1315e-01, -6.8645e-02, -2.1033e-01,  9.4513e-02,
         -7.9998e-02,  6.6883e-02,  5.2985e-02,  4.5739e-03,  1.0583e-01,
         -4.5220e-02, -9.0904e-03,  8.2827e-02, -1.3362e-01, -6.7235e-02,
          1.9438e-03, -4.3483e-02,  9.9083e-02, -3.4612e-02, -2.1234e-01,
          1.0221e-01, -9.0650e-02, -1.5209e-01, -9.4496e-02, -3.7238e-02,
         -1.1022e-01, -5.6732e-02,  3.5716e-02, -1.7685e-01,  9.0912e-02,
         -1.4253e-01, -1.0427e-02, -1.1439e-01, -6.9287e-02,  3.1953e-02,
         -1.4503e-01, -1.5553e-01, -1.8034e-01, -3.0496e-02, -1.0809e-02,
          1.2348e-01,  1.1634e-01,  1.7260e-01,  3.5692e-02, -4.9274e-02,
         -4.6776e-02, -1.4594e-01, -6.4116e-02,  5.4086e-02,  1.7549e-01,
         -1.7131e-01, -2.3566e-02,  1.3200e-01,  9.2775e-02,  2.8924e-02,
         -5.1050e-02,  4.4245e-02, -6.2847e-02,  3.1610e-02,  1.5044e-01,
          1.9344e-02, -7.9905e-02, -1.1045e-01,  1.7325e-01, -4.5421e-02,
         -1.3829e-01, -2.1175e-02,  2.4068e-01,  7.3709e-02, -1.1894e-01,
         -3.1301e-02,  1.0918e-01,  1.3093e-01,  7.9769e-02,  8.2108e-02,
          6.6651e-02,  3.0322e-02,  3.1324e-02,  7.4350e-02,  1.3370e-01,
         -1.1105e-01,  1.0952e-01,  1.6679e-02,  6.8369e-02,  5.1209e-03,
         -1.7720e-02, -1.0157e-01, -1.3004e-01,  6.1537e-02, -3.6965e-02,
         -5.5720e-03,  1.4211e-02, -3.3341e-02, -5.0988e-03,  3.5501e-02,
          1.1395e-01, -7.4218e-03, -1.2247e-01, -2.9845e-02,  3.3513e-02,
         -2.1570e-02, -4.8210e-02,  3.0376e-02, -6.4218e-02,  7.0922e-02,
          1.7718e-02, -6.8782e-02, -4.3030e-03,  7.0827e-02, -9.6241e-03,
          1.7542e-01, -2.0095e-02, -5.3108e-02,  1.5109e-01,  1.5682e-01,
          2.8846e-02, -4.6242e-02,  1.9079e-01, -2.0154e-02,  1.1266e-01,
          1.1151e-01, -1.2607e-01,  1.2059e-01,  4.5683e-02,  1.5597e-01,
         -3.6133e-02, -4.8355e-02,  5.5819e-02,  5.7645e-02, -4.0730e-02,
          1.4150e-01, -5.8886e-02, -1.5642e-01, -5.3169e-02, -9.6905e-02,
          1.3855e-01,  1.0479e-01, -3.7398e-02,  9.5933e-03,  1.3203e-01},
        '{-1.1491e-01,  9.8975e-03, -9.0949e-02,  9.0013e-02,  1.2665e-01,
         -1.6715e-01,  4.6048e-02,  4.7624e-02,  5.4970e-02, -1.0360e-01,
         -4.2058e-02, -2.0235e-02,  1.4650e-01,  1.0178e-01,  1.3315e-01,
          1.9568e-02,  8.9447e-02,  7.4470e-02,  5.8794e-02,  1.3796e-01,
         -2.6626e-01, -8.8388e-02, -7.9044e-02, -7.0410e-02, -2.0538e-02,
          6.6992e-02, -1.5414e-02, -5.6859e-02,  1.9764e-01, -2.4281e-02,
         -1.9080e-01, -4.2528e-01, -2.1985e-01,  2.9078e-03,  2.1740e-01,
         -1.3223e-02, -2.6241e-01, -3.4494e-02,  7.2087e-03, -1.6440e-02,
         -1.1968e-01,  4.2870e-02,  4.6711e-02, -1.9665e-02, -3.6315e-02,
          1.2818e-01, -5.5994e-02, -1.2628e-01, -9.1701e-02,  1.0578e-01,
          3.4534e-02,  4.5609e-03, -9.6287e-02, -2.8958e-02, -1.0803e-01,
          8.5483e-02,  9.6821e-02, -1.2095e-01, -1.3948e-01,  1.3421e-01,
         -8.7056e-02, -7.5676e-03,  4.8862e-02,  6.2714e-03,  2.1131e-01,
          1.7542e-01, -3.5177e-02,  3.4883e-02, -3.1952e-02,  1.6156e-01,
          6.2661e-02,  1.4136e-01,  1.0629e-01,  9.8876e-02,  4.6658e-02,
          6.5139e-02, -1.9882e-02,  5.2122e-02,  7.0502e-02,  2.7797e-01,
         -1.4804e-02,  4.5005e-02, -2.9799e-02,  1.2776e-01,  1.8865e-01,
          6.5252e-02,  1.6483e-01, -9.0665e-02,  7.3354e-02,  1.1429e-02,
         -4.4393e-02,  1.4427e-01,  2.1752e-02,  3.5977e-02, -8.7970e-02,
          4.2546e-02,  1.2797e-02,  7.6744e-03,  4.6300e-02, -9.0953e-02,
          1.1004e-01, -6.2268e-02,  1.1558e-01, -8.5039e-03,  1.2744e-01,
         -1.0172e-01,  6.5933e-02, -1.3608e-01, -1.8520e-01,  8.7010e-02,
          5.4846e-02,  1.4863e-01, -8.5294e-02, -7.5920e-03, -9.4880e-02,
          3.6291e-02,  9.4434e-02, -6.6694e-02,  1.3311e-01,  1.0720e-01,
         -1.0044e-01,  1.3860e-01,  1.9986e-02, -1.1085e-01, -1.0219e-01,
         -1.0719e-01, -2.0633e-01, -1.5040e-01, -7.6669e-02,  1.2631e-01,
         -1.3759e-01, -9.6417e-03, -8.9366e-02, -6.5166e-02,  3.8372e-02,
         -5.7268e-02,  1.5632e-02, -8.2192e-02,  8.9298e-03,  1.4205e-03,
          1.1881e-01, -1.0502e-01,  6.5675e-02,  4.1302e-02,  1.6545e-01,
         -8.9264e-02,  9.7108e-03,  5.2869e-02,  3.2239e-02, -2.3433e-02,
          3.2842e-02,  8.4551e-02,  1.2771e-01,  9.3593e-03,  7.1677e-02,
         -4.9618e-02,  1.8004e-01,  7.2197e-06, -1.9865e-03, -1.2002e-01,
          1.1905e-02, -7.7872e-04, -9.3492e-02, -1.3362e-01,  1.0904e-01,
          1.4168e-01,  1.6880e-01,  5.9445e-02,  1.6384e-01, -9.8388e-02,
          7.3235e-02,  5.9703e-02,  1.7063e-02,  1.6037e-01, -4.4810e-02,
         -9.0209e-02, -6.6820e-02, -1.4584e-01, -3.4877e-02,  2.2178e-02,
          6.9512e-02, -4.0707e-02,  1.0277e-01,  3.4602e-02, -9.9834e-02,
          1.4957e-01,  1.8641e-01, -3.6456e-02, -1.6503e-01,  6.6795e-02,
          2.5145e-02,  1.6652e-01, -1.8074e-02, -8.6670e-02, -9.3954e-02,
         -8.6859e-02, -7.3930e-02,  1.1867e-01,  8.8946e-03, -1.0645e-01},
        '{-5.1013e-02, -5.1930e-02, -6.7805e-02,  1.7860e-02, -1.4975e-01,
          8.9135e-02,  1.5433e-01,  9.4606e-02, -1.2199e-02,  1.2962e-01,
         -3.3248e-03,  5.1932e-02,  1.0756e-02,  9.9867e-02, -1.0868e-01,
          8.9914e-02,  1.0561e-01, -5.1985e-02, -9.9533e-02, -5.8649e-02,
          3.4227e-03, -7.7476e-02,  2.7341e-02,  4.7153e-02, -3.4749e-02,
         -2.3581e-02, -3.5644e-02,  3.2702e-02,  8.1514e-02,  1.2221e-01,
          1.5871e-02,  3.0017e-02,  9.9218e-02,  8.5806e-02,  4.5630e-02,
         -2.4328e-02, -7.1619e-02, -8.4650e-02,  6.2320e-03,  9.3056e-02,
          3.9883e-02,  1.0438e-02,  1.0380e-01, -1.0861e-01, -9.8768e-02,
          8.5543e-02, -2.6775e-02, -2.1049e-02, -9.1751e-02,  1.3264e-02,
          3.8827e-02,  7.3867e-03, -1.6029e-01, -1.2846e-01, -9.3388e-02,
          9.7360e-02,  3.2489e-02,  2.1381e-02, -1.3631e-02, -2.2709e-02,
          7.5750e-02,  3.9726e-02,  5.9075e-02, -7.1155e-02,  1.1347e-01,
         -5.7139e-02,  6.3272e-03,  5.9542e-04,  4.4412e-02, -3.1660e-03,
         -8.0316e-02,  3.2092e-02,  5.8564e-02, -1.7102e-03,  4.4561e-02,
          2.7660e-02,  2.3260e-02, -9.9845e-02, -1.3491e-01, -8.1259e-02,
          1.3983e-02,  3.0600e-02, -1.2868e-01, -1.1009e-01, -4.2556e-02,
          1.0702e-02,  6.1267e-02, -1.0648e-02, -5.4690e-02, -4.9519e-02,
          3.5894e-02,  5.6010e-02, -6.7543e-02,  2.5094e-02,  9.0557e-02,
         -2.8447e-02, -4.3920e-03,  9.2484e-03,  7.7130e-02,  7.4364e-02,
          3.4056e-03,  5.3668e-02,  5.5494e-02, -1.2693e-01,  5.1120e-02,
         -6.6875e-02,  9.4124e-02, -2.8082e-02,  4.2366e-02, -1.7277e-02,
          3.9165e-02,  1.0797e-01,  5.6388e-03, -1.5540e-04, -1.5986e-02,
         -1.8903e-02,  1.3995e-01, -2.9178e-02, -7.2442e-02, -1.0980e-01,
          2.7613e-03, -1.9391e-02, -7.9176e-03, -2.4119e-02,  1.4624e-01,
         -2.6080e-03,  2.8247e-03,  1.8717e-02,  5.1081e-02,  4.4505e-02,
          4.7523e-02,  5.4782e-02, -1.5547e-03,  9.3718e-03,  2.7851e-02,
         -3.2341e-02, -2.2786e-04, -3.3611e-02,  3.8710e-02,  3.3884e-02,
          5.4010e-02,  5.2369e-02, -9.0819e-04,  8.1491e-03, -4.3164e-03,
         -1.6898e-02,  1.1486e-02, -3.3261e-02, -2.2903e-02, -7.5603e-03,
         -8.5795e-02,  8.7261e-02, -3.9834e-02, -7.5157e-02, -1.2931e-01,
         -7.7337e-02, -8.9414e-03, -2.4927e-02,  1.5381e-02,  1.1775e-03,
         -1.3930e-02,  5.1246e-02, -9.6348e-02, -4.7431e-02, -1.1263e-01,
          6.1470e-02,  1.4684e-01, -1.0359e-01, -1.2835e-01,  1.0618e-01,
          1.2075e-02, -5.3314e-02, -5.0075e-03, -4.5303e-02, -1.5839e-02,
          8.0957e-02, -3.8532e-02,  9.8745e-03,  1.9714e-02, -5.5501e-02,
          1.2278e-01,  3.3439e-02, -3.3542e-02, -5.7444e-02,  9.6559e-02,
         -6.8967e-03,  4.8349e-02, -5.1472e-03,  2.3489e-02,  7.5612e-02,
         -1.1173e-01, -2.4169e-04,  7.2070e-02,  3.1593e-02,  1.1870e-01,
         -5.3013e-02, -6.7265e-02,  6.6470e-02, -8.3994e-02,  1.4755e-01},
        '{-8.2088e-02,  1.0307e-01, -9.0172e-02, -4.1279e-02,  1.3074e-01,
          9.2532e-02, -2.5678e-02,  1.2066e-01,  2.1909e-01, -1.1227e-01,
         -6.0523e-02, -1.3452e-01, -1.1416e-01,  1.9077e-02, -2.1976e-01,
          1.4716e-01, -1.2038e-01,  2.2911e-02,  1.0566e-01, -7.8994e-02,
         -1.3579e-01, -1.2114e-02,  1.0250e-01, -9.6476e-02,  1.7883e-01,
          1.9708e-01,  1.9514e-01,  9.4386e-02,  3.4774e-02, -2.5080e-01,
          3.2562e-03,  2.9097e-02,  2.6125e-01,  5.3973e-02, -2.8379e-01,
          1.1521e-01,  2.3179e-01,  1.4619e-01, -2.5910e-03, -9.9177e-02,
         -1.8149e-02,  4.0842e-02, -4.4901e-02,  7.0621e-02,  6.6392e-02,
          7.5349e-02, -2.0798e-01,  1.8777e-02, -7.9810e-03,  1.8924e-02,
         -1.9170e-02,  1.9537e-03, -2.0800e-03,  2.0627e-02, -9.4994e-03,
         -8.4327e-02,  1.5023e-02,  6.2521e-02,  9.1471e-02,  8.9047e-02,
         -1.6417e-02,  9.3950e-02, -2.7156e-02,  1.4228e-02,  1.5840e-02,
          4.0174e-02,  7.1398e-02, -1.7997e-01, -2.3556e-01, -5.3242e-02,
         -1.3471e-01, -3.9721e-02, -1.0597e-01,  1.2105e-01,  1.6816e-01,
          1.5001e-02, -2.1665e-02, -1.2867e-01,  5.3222e-02, -8.1387e-02,
         -7.5112e-02, -1.4634e-01, -2.8978e-02,  8.5847e-02, -9.4423e-03,
         -7.2836e-03, -1.4701e-01,  8.2263e-02,  1.3524e-02,  1.0542e-01,
         -3.0934e-02,  6.3359e-02,  8.4343e-02,  4.4300e-02,  5.5630e-03,
         -7.0018e-02,  3.0439e-02, -1.0217e-01,  1.4535e-02, -9.5770e-03,
         -1.2150e-01, -1.5491e-02, -4.4370e-03,  1.1098e-01, -1.0834e-01,
          5.3259e-02,  3.4864e-02,  1.3680e-01,  1.5421e-01,  1.7393e-01,
          5.8354e-02, -1.8918e-01, -7.5100e-02,  1.7294e-01,  1.3294e-01,
         -9.2310e-02,  5.4436e-02,  2.2045e-03,  1.5547e-01, -1.5944e-01,
          7.8005e-02, -9.3053e-02,  1.0928e-02,  5.7126e-02, -8.5112e-02,
          1.2521e-01,  5.4675e-02,  1.3544e-01,  6.1565e-02, -1.2855e-01,
         -3.3227e-02,  1.7759e-01,  1.1256e-01,  2.1084e-01, -5.0122e-02,
          1.8904e-01,  1.1723e-01, -8.3622e-02,  6.1367e-02,  8.3065e-02,
         -1.4592e-01,  1.6460e-02, -1.6459e-01,  1.0738e-01,  2.6352e-02,
         -1.6136e-01, -7.6032e-02, -4.2221e-02, -9.9027e-02, -3.8263e-02,
          1.7694e-02,  1.1886e-01,  1.2374e-01,  1.5581e-02, -3.4067e-02,
          1.0864e-01, -7.3345e-02, -6.5148e-02,  1.2140e-01, -8.4215e-02,
         -5.8847e-02, -2.6603e-02,  3.8992e-02,  4.8207e-02,  3.9285e-02,
         -7.4956e-02, -4.1747e-02,  1.2425e-01,  4.6243e-02, -4.9955e-02,
          9.1594e-02,  1.0928e-01,  4.1429e-02, -8.2226e-02, -6.1136e-02,
         -2.4292e-03, -9.0924e-02,  6.2366e-02, -1.6290e-02, -5.1476e-02,
         -1.2840e-01, -3.5174e-02,  1.5429e-02, -3.7443e-02,  1.7409e-01,
          2.2433e-02, -3.6753e-02,  1.5569e-03, -9.1048e-02,  5.1168e-03,
          3.1571e-02,  2.7241e-02,  1.5809e-01,  9.7499e-02, -1.4902e-02,
          1.2081e-02, -1.2581e-01,  1.1178e-01, -3.3755e-02,  3.7831e-02},
        '{ 5.7475e-02,  1.0813e-01,  2.2457e-02,  3.8585e-02,  1.9115e-01,
          1.3240e-01,  2.3650e-02, -3.2054e-02, -1.4510e-02,  1.9655e-02,
         -2.0674e-02,  4.4006e-02, -8.3206e-02, -1.3403e-01,  1.1134e-01,
          2.0484e-02, -1.5012e-01, -1.1536e-01, -4.5246e-02,  5.7024e-03,
         -5.7547e-02, -4.8497e-02,  1.1679e-01,  1.5918e-02, -1.4253e-01,
          5.5990e-02,  1.0095e-01, -1.1996e-01, -7.7799e-02, -3.2153e-01,
          3.4473e-02,  1.1968e-02, -1.1236e-02, -1.4455e-01, -3.2977e-01,
          3.3342e-03, -1.7597e-01, -1.4330e-01, -7.2610e-02,  7.5424e-02,
          6.5078e-02,  2.9216e-02, -7.6860e-02,  2.0866e-02, -1.5291e-02,
         -1.3939e-01, -6.2201e-02, -9.2871e-02, -1.3152e-01, -1.0748e-01,
         -1.4349e-01, -1.3700e-01,  8.3992e-02,  3.7452e-02, -8.5764e-03,
          1.3286e-01,  1.6729e-01, -5.4063e-02,  1.1070e-01, -1.6300e-01,
          7.3220e-02,  2.2456e-02,  9.3360e-02,  9.2803e-02,  4.8044e-02,
          1.4376e-01, -7.7416e-02,  6.5673e-02,  1.0077e-01,  7.9328e-02,
         -1.1510e-02, -1.2810e-02,  2.4403e-02, -9.7729e-02,  2.1426e-02,
         -1.3778e-02, -5.5860e-02,  2.1129e-04, -3.5434e-02,  4.7107e-02,
          5.3457e-02,  3.6826e-02,  1.1382e-01, -2.3152e-03,  1.1228e-01,
         -8.6915e-02, -9.7274e-02, -7.8199e-02,  4.3965e-02,  1.3382e-02,
          1.6604e-02,  1.0933e-01, -2.7368e-02,  4.3144e-02, -1.2153e-01,
          9.3698e-03,  4.4583e-02,  8.1610e-02,  1.5429e-02,  9.4815e-02,
          9.7081e-02, -7.0907e-02, -5.7389e-02, -1.0836e-01,  1.7972e-01,
         -2.9774e-02,  8.2993e-02,  7.4138e-03,  1.1846e-01,  3.9896e-02,
          1.5456e-01,  1.6626e-01,  1.6226e-01, -1.8445e-03,  8.5288e-02,
          1.7720e-01,  5.1412e-03, -1.4094e-02, -7.0793e-02, -9.8426e-02,
         -1.0978e-01,  1.1286e-01,  6.2787e-02,  1.3583e-01,  1.6597e-02,
         -1.7111e-01, -1.3504e-01, -1.5232e-02, -6.6112e-02, -8.0615e-02,
          2.9100e-02,  2.5575e-02, -1.2650e-01,  6.5780e-02, -6.8634e-02,
         -2.5360e-02,  1.3416e-01, -9.8206e-02,  5.1954e-02,  1.2257e-01,
          6.4431e-02,  1.3085e-01, -2.5931e-02,  1.0942e-01, -7.2406e-03,
          7.9495e-02, -1.0579e-01, -1.3669e-01, -3.3778e-02, -6.7862e-02,
          4.5548e-02,  1.5729e-01,  3.9734e-02,  1.5296e-01,  6.8285e-03,
          9.4934e-02,  1.5201e-01,  4.7953e-02, -9.2203e-02,  1.3169e-01,
         -9.0950e-02,  1.0137e-01, -7.6983e-02, -5.0561e-02, -5.7249e-02,
          5.6278e-02, -6.8416e-02, -8.5421e-02,  1.9942e-03,  5.9096e-02,
         -6.6719e-02, -9.3265e-02, -7.6698e-02, -2.8109e-02,  4.6492e-03,
         -3.8130e-02,  1.5555e-01,  9.7290e-02, -1.0410e-01, -7.4924e-03,
          1.0612e-01, -1.2947e-01, -6.0895e-02,  1.0459e-01, -4.2177e-02,
         -8.4109e-02, -1.1365e-01, -1.5917e-02, -3.1450e-02,  1.1360e-01,
          3.8720e-02,  8.2997e-02, -6.2159e-02,  1.1974e-01,  5.1319e-02,
         -8.7519e-02, -1.2608e-01, -1.3557e-01,  1.1001e-01, -1.1529e-01},
        '{ 1.2991e-01, -1.1682e-01, -7.9969e-02,  1.1858e-01, -9.7086e-02,
         -1.3317e-01,  1.1238e-01, -7.9846e-02,  8.5076e-02,  1.5891e-02,
          1.1384e-01,  9.1233e-02,  1.0854e-01,  1.3442e-01,  1.6496e-01,
          1.3669e-01,  1.7991e-01,  1.7892e-01, -7.2141e-02, -8.0940e-02,
         -4.7053e-02, -2.0557e-02, -4.4221e-02, -1.1258e-02,  6.0256e-02,
         -2.6475e-02,  1.6584e-01, -9.1156e-02,  1.6627e-02,  1.7305e-01,
         -1.1658e-01, -3.5535e-02,  2.1129e-01,  5.1471e-02,  1.3017e-01,
         -1.7690e-01,  7.3635e-02, -1.2578e-01,  2.9550e-02, -9.9510e-02,
         -1.5404e-02,  7.0993e-02,  1.3061e-01, -1.5330e-01, -1.1432e-01,
          1.1481e-01,  2.6688e-01,  1.9642e-01,  1.2732e-01, -1.4668e-02,
         -1.4016e-01, -3.6546e-02, -9.0454e-02, -6.2611e-02, -7.1859e-02,
         -1.2983e-01, -6.8087e-02,  3.7106e-02,  9.7595e-02,  9.1178e-02,
          4.8506e-02,  9.2337e-02, -1.9944e-02,  2.0028e-01,  1.8944e-02,
          2.3326e-02, -8.8291e-02,  1.4320e-01,  2.9508e-02,  2.7177e-02,
          5.6403e-02,  2.6201e-02,  7.7019e-02, -5.6722e-02,  8.9848e-02,
         -3.8650e-02, -1.4061e-01, -7.7478e-02, -1.5703e-01, -4.8556e-02,
          4.3218e-02,  1.3600e-01,  1.4631e-02, -8.6596e-02, -1.9248e-01,
          1.6929e-04,  1.2617e-01, -1.0558e-02, -7.4792e-02, -1.8370e-03,
         -1.4318e-01, -5.3878e-02, -9.8794e-02,  5.1445e-02, -4.3922e-04,
         -1.4598e-01, -3.8430e-02, -1.0168e-01,  4.1060e-02, -6.6876e-02,
         -1.4157e-01,  6.2679e-02, -4.9551e-02,  4.3822e-02, -1.5608e-02,
         -1.2007e-01,  1.2898e-01, -1.2878e-01,  3.4858e-02, -7.4571e-02,
         -2.2074e-02,  1.3171e-01, -1.5247e-01, -8.4275e-02,  4.7467e-02,
         -9.4087e-02,  9.1211e-02, -7.9593e-02,  2.3827e-02,  1.8135e-01,
          1.8433e-02,  5.5026e-02, -1.0425e-02, -5.3994e-02, -7.5748e-03,
         -9.5260e-02, -8.7474e-02,  1.0078e-01,  1.2709e-01,  2.6712e-02,
          3.7861e-02,  9.0025e-03, -1.2796e-01,  1.4333e-01, -6.2511e-02,
         -5.1823e-02,  3.7837e-02,  3.6748e-02,  1.1024e-01, -1.0972e-02,
          9.6672e-02,  1.7995e-01,  1.0262e-01, -2.0913e-02,  6.1980e-02,
          1.0407e-01,  8.6942e-02, -2.7034e-02,  1.0454e-01,  6.7402e-03,
         -1.4330e-01,  7.8993e-02, -1.7362e-02,  1.1680e-01, -1.9867e-02,
          9.6848e-02,  1.2099e-01, -5.5024e-02,  2.7299e-02, -7.3496e-02,
         -9.2674e-02,  9.6538e-02,  1.0679e-01,  6.8710e-02,  4.0637e-02,
          2.3044e-02, -5.3897e-02, -1.1973e-01, -2.6723e-02, -8.3382e-02,
          6.1312e-02,  1.6678e-01,  7.4251e-02,  1.6005e-03,  1.0839e-01,
          9.9324e-02,  1.0335e-01,  1.8058e-01,  4.0409e-03,  6.4109e-02,
          1.2191e-03, -9.6053e-02, -1.2070e-01, -4.0487e-02,  1.4945e-01,
          1.1471e-01, -4.7097e-02,  7.1803e-02, -5.0058e-02,  9.7168e-02,
         -6.1393e-02,  5.0080e-03,  2.7569e-02, -3.3845e-02,  1.0782e-01,
          5.8593e-02, -9.9623e-02, -1.2157e-02, -7.0098e-02, -3.6889e-02},
        '{ 9.5079e-05, -7.7471e-02, -1.2349e-01, -2.3192e-02,  1.0399e-01,
         -7.4014e-02, -3.3031e-02, -8.3854e-02,  5.9693e-03, -6.6467e-02,
          7.4103e-03,  1.1234e-01,  8.0723e-02,  1.0941e-01, -1.6680e-03,
          1.6338e-01,  1.1240e-01,  1.6516e-01,  1.1789e-01, -3.8583e-03,
         -8.5879e-02,  9.6700e-02,  1.2113e-01,  1.5617e-01,  2.4750e-01,
          1.4407e-01,  5.0104e-02, -5.7261e-02,  1.6001e-01,  2.8435e-01,
         -2.4557e-01, -5.6062e-02, -1.3271e-01,  2.7171e-01,  3.4082e-01,
          1.9100e-01, -4.7906e-02, -2.2817e-02,  4.2057e-02,  2.7568e-01,
          1.1475e-01, -2.6229e-01,  2.8032e-03,  4.8714e-03, -2.9314e-01,
         -9.7545e-02,  1.1324e-01, -1.3030e-01, -1.6686e-01, -1.1399e-01,
          5.6408e-02, -4.4058e-02, -5.2068e-02, -8.1566e-02, -1.5225e-01,
          1.6665e-01,  4.2327e-02,  1.5314e-01, -1.8773e-01,  8.9949e-02,
          1.4269e-01,  1.4918e-01,  7.3914e-02, -2.0295e-01,  3.1413e-01,
          1.1403e-01,  3.3196e-02,  7.4195e-02,  1.4726e-01, -1.5846e-02,
          1.6066e-01,  1.0004e-01, -2.1462e-02,  1.4489e-01, -6.4337e-02,
          1.9631e-02,  6.2070e-02,  6.3688e-02,  6.8973e-02, -5.0656e-02,
          1.5228e-01,  9.2093e-02, -5.0453e-02, -1.0109e-01, -1.9773e-01,
          9.7407e-02, -2.9783e-02,  9.2791e-02, -2.1375e-01, -1.1909e-01,
          1.6944e-03, -7.4702e-02,  3.0509e-02, -1.0246e-01,  1.2215e-02,
          1.2519e-01,  1.2074e-01, -9.2300e-02,  1.1859e-02,  1.0432e-01,
         -9.8452e-02,  5.1492e-02,  2.0991e-01,  8.9301e-02,  7.4948e-02,
          5.1653e-02, -1.0148e-01,  1.4206e-01,  3.7801e-02,  2.5313e-02,
          2.2673e-02,  1.0124e-01,  1.0512e-01,  8.9701e-02, -8.1039e-02,
         -6.9977e-02,  6.5663e-02, -3.5362e-02, -1.2470e-01,  6.6675e-02,
         -6.4484e-02,  6.4122e-02,  2.6366e-02,  2.1021e-01,  1.3518e-01,
          4.9662e-02,  3.4717e-02,  7.1074e-02,  1.0125e-01,  3.1181e-01,
          4.2473e-02, -7.4685e-02, -8.5167e-02,  7.2001e-02,  1.2360e-01,
         -5.9321e-02,  7.8402e-02,  7.5614e-02,  1.1591e-02,  1.3290e-01,
          1.1613e-02, -1.2097e-01, -1.2147e-02,  5.6642e-02, -1.3565e-01,
          1.0783e-01,  1.9067e-01,  7.5245e-02,  1.2553e-01,  2.1360e-03,
          5.2046e-02,  5.0204e-02,  2.2181e-01, -2.2981e-02, -6.2953e-02,
          5.5409e-02, -1.4895e-01, -7.1490e-02, -9.3964e-02,  1.3228e-02,
         -1.6377e-01,  3.7466e-02,  1.1818e-01, -9.7402e-02, -3.0027e-02,
         -6.3026e-02,  8.6706e-02, -8.3204e-02,  8.7320e-02, -7.8349e-02,
          1.4875e-01,  1.6507e-01,  1.6978e-01,  1.0524e-01,  2.5765e-01,
         -1.5349e-01,  1.6805e-01,  4.3581e-04, -2.7541e-02,  1.6948e-01,
         -5.4085e-03, -1.4298e-01, -5.2654e-02, -3.2834e-02, -5.3137e-03,
         -1.3690e-01,  1.0751e-02,  8.0819e-02, -1.2759e-02, -1.4254e-01,
         -1.6456e-01, -4.8748e-02,  8.6785e-02, -7.1214e-03,  8.2884e-02,
          1.2404e-01,  1.6201e-01,  4.2853e-02, -1.7054e-02, -2.0336e-02},
        '{-1.7137e-01, -5.7594e-02,  1.8437e-01,  1.0537e-01,  5.8545e-02,
          9.2523e-03, -5.8363e-02,  3.5234e-02,  6.9971e-02,  1.4287e-01,
          1.0047e-01,  2.2854e-02,  1.6223e-01, -7.3317e-02, -9.9027e-02,
          1.4393e-02, -7.1785e-02,  5.7721e-02, -2.5191e-02,  4.8604e-04,
         -1.7544e-02,  2.4485e-02, -5.4031e-02, -6.6292e-02,  2.3380e-01,
          7.9135e-02,  1.2213e-01, -1.3513e-01, -1.3139e-01, -3.8053e-03,
          9.9060e-02, -1.9222e-01,  5.8078e-02, -4.2081e-02, -6.9666e-02,
          7.4370e-02,  1.2001e-01, -1.9476e-01, -5.7709e-02, -1.1054e-01,
         -3.0763e-02, -3.1201e-01, -7.3818e-02,  8.5167e-02,  9.9087e-02,
         -1.2233e-03, -4.9366e-02, -1.6536e-01, -8.5963e-02, -1.1717e-02,
         -4.1971e-02, -7.3333e-02,  1.3179e-01,  9.3103e-02,  5.8456e-02,
         -1.1104e-01, -4.3943e-02,  4.7644e-02,  5.9248e-02,  1.5029e-01,
          1.5053e-01, -3.7861e-02,  9.2767e-02, -4.8766e-02,  4.2529e-02,
          5.6006e-02, -1.1651e-01, -8.2312e-02,  6.6293e-03,  5.7730e-02,
          4.3381e-02,  5.2548e-02, -1.3520e-01,  1.2214e-01,  8.2782e-02,
          8.7813e-02, -1.0653e-03,  1.3016e-01, -1.0908e-01, -1.6774e-01,
         -1.1260e-01,  1.1278e-01, -1.0615e-01,  3.8022e-03,  7.1504e-03,
          1.2989e-01, -1.1863e-01, -3.6552e-02,  6.5279e-02,  2.4658e-01,
          1.7375e-02, -3.5538e-02,  3.7585e-02, -3.8700e-04,  1.1180e-01,
          4.4804e-02,  1.7651e-02, -2.8888e-02, -2.0283e-02,  7.8417e-02,
         -1.3367e-01,  6.1273e-02, -6.6736e-02, -4.3296e-02,  1.7495e-01,
          1.0413e-01,  9.9697e-02,  3.9223e-02,  9.8603e-02,  1.4992e-01,
          4.2078e-02,  1.3056e-01,  2.5862e-02, -8.1303e-02,  1.2382e-01,
         -2.2596e-02,  1.4617e-01,  1.4651e-01,  4.1308e-02, -3.7950e-02,
          1.4797e-01,  1.7021e-01,  9.1621e-02,  9.2418e-03,  1.6737e-01,
         -6.9543e-02, -3.5446e-02,  1.6225e-01,  2.6909e-02,  2.7636e-03,
          5.6546e-02,  4.3033e-02, -1.4871e-03,  1.0420e-01, -1.6651e-01,
          1.0189e-01, -1.0261e-01, -1.4394e-01, -5.4484e-02,  4.9146e-02,
         -1.7927e-01, -8.3510e-03, -5.6117e-02,  3.7649e-02, -2.1635e-02,
          2.7333e-02,  6.1627e-03, -1.4170e-01, -1.6236e-01,  1.2924e-01,
          4.9066e-02, -8.1253e-03,  4.4207e-02,  1.8039e-04, -8.7672e-02,
          4.5629e-02, -1.1149e-01, -5.7776e-02, -1.4391e-01,  8.5333e-02,
          8.1024e-02,  1.1185e-01, -6.9760e-02, -1.1328e-01, -6.4369e-02,
         -4.4665e-02,  1.8436e-01,  1.3284e-01,  9.3340e-02, -6.1283e-02,
         -3.3195e-02,  9.7008e-02,  7.0031e-02, -7.3381e-02,  9.6421e-02,
         -6.1443e-03, -1.3188e-01, -7.5016e-02, -5.7621e-02, -3.8031e-02,
         -4.5560e-02,  9.4655e-02, -1.1421e-01,  2.8390e-02, -3.6281e-02,
          5.7355e-02, -8.5650e-02, -8.6325e-02, -1.2488e-01, -4.5025e-03,
         -8.1771e-02,  1.6414e-01,  3.7653e-02, -5.3373e-02,  4.5397e-02,
          1.3818e-01,  7.7858e-02,  6.9618e-02, -6.0317e-02, -5.4634e-02},
        '{-1.4806e-01, -1.6292e-02, -8.9363e-02,  5.9800e-02,  5.1147e-02,
          2.3799e-02,  1.2969e-01, -8.2215e-02, -1.1910e-01, -1.0354e-01,
         -3.9366e-02, -5.8611e-02, -6.8580e-02,  1.2727e-01, -4.5116e-02,
         -4.5057e-02,  1.3935e-02, -3.6901e-02, -1.2338e-01, -5.6898e-02,
         -1.2003e-02,  1.5889e-01,  1.6371e-01, -7.0386e-02,  1.4190e-01,
         -2.3525e-02, -1.3694e-01,  4.9913e-02,  2.8788e-01,  2.7132e-01,
         -1.9178e-01, -1.4169e-01,  6.7468e-02,  8.5683e-02,  2.6975e-01,
         -1.8925e-01, -2.0868e-01,  6.7502e-02,  1.6733e-02,  8.6424e-02,
          8.9442e-02,  1.2695e-01, -4.4275e-02,  4.9647e-02, -1.6227e-01,
          7.6027e-02,  2.7905e-02,  2.2227e-01,  1.9706e-01, -4.2111e-04,
          2.2417e-02,  9.0102e-02,  1.0166e-01, -1.5526e-01, -3.8946e-02,
         -1.0956e-01,  3.0051e-02,  2.1971e-02, -5.2516e-02, -2.2678e-02,
         -1.0048e-01,  1.0791e-01, -8.4057e-02, -2.7803e-02,  1.3291e-01,
         -6.8774e-02,  9.9523e-02, -1.0271e-01, -2.4755e-02,  1.0700e-02,
         -1.0250e-01, -1.8187e-02, -1.4336e-02, -3.6539e-02,  6.8373e-02,
          2.7054e-02, -4.8509e-02,  1.7199e-02,  1.2924e-01,  6.9518e-02,
          3.9517e-02,  7.7369e-02,  5.9804e-02, -4.1500e-02,  1.9710e-02,
         -6.2825e-02,  6.8959e-02, -9.8927e-03, -9.7492e-03, -1.9901e-01,
         -9.0203e-02,  8.8761e-03, -1.2614e-02,  1.5875e-01,  1.6188e-01,
         -1.3000e-01, -2.9460e-02,  1.8198e-02,  5.7737e-02, -1.2746e-02,
         -3.2292e-02,  2.1179e-02,  4.3251e-03, -9.5506e-02,  2.1887e-04,
         -1.4013e-01, -6.5425e-03,  3.8628e-02, -1.2873e-01,  1.0740e-01,
          1.4029e-01,  2.6238e-02,  6.4422e-02, -1.4177e-01,  5.6621e-04,
          1.1110e-01,  2.1819e-03,  2.9086e-02, -8.2813e-02, -1.0786e-01,
          3.2675e-02,  5.1494e-02,  1.2948e-01,  1.6147e-01,  8.2937e-03,
          1.1822e-01,  4.1296e-02, -1.0185e-01,  1.1516e-01,  1.3840e-04,
         -1.9010e-01, -2.4854e-02, -8.7637e-03, -7.8581e-05,  1.5537e-01,
         -2.8270e-02, -8.4795e-03,  5.7166e-03,  4.8199e-02,  4.4708e-03,
          3.2541e-02,  4.4041e-02, -6.9758e-02,  4.6798e-02,  8.7750e-03,
          1.1450e-01,  3.9567e-02,  7.0607e-02, -5.6345e-02,  1.9559e-02,
         -2.8957e-02,  1.6733e-02,  8.0252e-02, -9.8545e-02,  8.8639e-02,
          2.5568e-02, -6.3340e-03,  1.7894e-01,  4.8239e-02, -9.2657e-02,
          1.0926e-01, -7.4840e-02, -1.2879e-01, -1.4566e-01,  7.2032e-03,
         -2.0082e-03, -6.4236e-02, -1.7180e-01, -8.7875e-02, -6.5859e-02,
          7.4770e-03, -2.2577e-02,  1.1619e-01,  6.8593e-02,  1.7499e-01,
          6.5894e-02,  8.7992e-02,  8.1183e-02, -3.0097e-02,  9.6706e-02,
          4.3289e-02, -1.3961e-02,  8.4332e-02, -1.8170e-02, -9.0314e-02,
         -2.6531e-03,  1.7070e-01,  3.0044e-02, -1.0159e-01,  3.3763e-02,
         -8.3898e-03,  1.1880e-01, -3.7295e-02, -1.1497e-01, -3.7958e-02,
         -6.0090e-02, -3.6203e-02, -3.3091e-02,  1.1259e-01, -2.1728e-03},
        '{-9.2445e-02, -1.3900e-01, -1.2760e-01,  9.2934e-02, -4.3527e-02,
          6.1342e-02,  2.2067e-02, -3.2714e-02,  6.8051e-02,  3.3231e-02,
          1.9224e-01,  1.2371e-01, -4.9558e-02,  4.6393e-02,  6.9602e-02,
          5.9058e-02, -1.0036e-01,  4.3626e-02, -4.2402e-02,  3.2073e-02,
          6.0017e-02, -9.4827e-02, -1.2811e-01, -1.5848e-01, -1.3425e-01,
          1.5922e-01,  1.0614e-01,  3.4813e-02, -2.1084e-02, -6.4171e-02,
          1.9168e-01, -5.9602e-02,  9.0000e-02,  3.8349e-03, -2.1803e-01,
         -4.7810e-02,  4.8444e-02,  8.0143e-02, -1.5479e-01, -1.1903e-01,
         -2.3702e-02,  2.2010e-01,  8.9044e-02,  7.2159e-02,  2.4329e-01,
         -8.6172e-02,  1.0908e-01,  2.3380e-03,  1.8999e-01,  1.1254e-01,
         -4.5437e-02, -1.5625e-02, -4.6330e-02,  1.1236e-01, -3.6876e-02,
         -4.7434e-02, -2.1196e-02,  1.2383e-01,  1.1413e-02, -5.9349e-03,
         -8.3905e-02,  5.2644e-03,  1.6210e-02,  1.7346e-02, -1.9462e-01,
         -7.8732e-02,  2.4534e-02,  1.4645e-01,  7.7537e-02,  1.0229e-01,
         -5.8788e-02, -2.2841e-02, -3.5052e-02, -4.5906e-03,  1.6760e-01,
          1.5066e-02, -1.3573e-01, -2.3444e-02, -9.6094e-02,  1.0449e-01,
         -6.1384e-02, -7.1670e-02, -3.1206e-02,  2.7470e-02,  4.2878e-02,
          8.2954e-02, -1.4664e-02, -8.3478e-02,  8.0342e-02,  1.0044e-01,
          1.4667e-01,  3.9651e-02,  4.7227e-03,  7.1278e-02,  2.6273e-02,
          9.7702e-03, -6.1449e-02,  7.8525e-02,  1.6666e-02, -2.2047e-01,
         -1.6395e-02,  2.0261e-02, -1.2684e-01, -5.7320e-02, -4.1932e-02,
         -1.6412e-02, -1.0911e-01,  6.3510e-02, -4.3059e-02, -6.2393e-02,
         -6.5037e-02,  8.7975e-02, -7.3036e-02, -2.5111e-02, -3.9560e-02,
         -1.1247e-02,  1.4914e-02,  1.2104e-01,  9.9765e-03, -2.2015e-02,
          2.7573e-02, -2.7933e-02, -8.1685e-02, -4.2664e-02,  3.1008e-02,
         -5.2608e-02,  4.0470e-03,  1.2349e-02, -1.9140e-02, -1.0841e-01,
          3.6728e-02,  1.3165e-02, -3.1675e-02, -4.5682e-02,  2.5177e-02,
         -1.6617e-01, -3.1123e-03, -4.4712e-04,  4.4629e-02, -1.5514e-01,
          6.1462e-02,  8.0443e-02, -4.6083e-02,  2.8830e-02,  6.4720e-02,
         -1.1671e-02, -3.1214e-02,  2.7049e-02,  3.9839e-02, -4.7468e-02,
         -3.2234e-02, -8.2680e-02,  5.1808e-02, -9.0132e-02,  2.9700e-02,
         -6.2253e-02, -8.5063e-03,  8.4091e-02,  7.5523e-02, -8.4452e-02,
          1.2309e-01,  1.0751e-01,  1.5746e-01, -5.6412e-02,  6.4483e-02,
         -3.9681e-02,  8.2830e-02, -8.7541e-02,  1.1040e-01,  1.0286e-01,
         -7.5159e-03, -1.1361e-01,  5.2102e-02,  3.8387e-02, -1.4000e-01,
          2.2090e-02, -7.9218e-03,  3.7081e-02, -8.4697e-02, -5.2771e-02,
         -3.1912e-02, -9.5795e-02, -7.5231e-02, -1.0149e-01, -1.5845e-01,
          7.0459e-02,  1.8174e-01,  1.5917e-01,  1.3563e-01, -1.0017e-01,
         -3.1921e-02,  4.9870e-02,  8.4621e-02, -6.1998e-02,  7.7268e-02,
         -1.2704e-01,  6.4057e-02, -7.3533e-02,  7.3043e-03, -1.4329e-01},
        '{-1.9232e-01,  4.7268e-02,  6.0244e-02,  1.8697e-01, -3.1384e-02,
          6.9528e-02,  1.5623e-01, -1.3450e-01, -1.0634e-01,  1.0138e-01,
         -1.1420e-01,  1.2244e-02, -6.7737e-02, -8.0989e-02, -5.1501e-02,
         -2.8023e-01, -4.9008e-02, -1.2772e-01, -7.5640e-02, -1.0601e-02,
         -3.4483e-02, -2.1942e-01, -5.5893e-02, -2.9476e-02,  6.9061e-03,
         -1.1144e-01, -1.0082e-01, -2.4232e-01, -2.3663e-01,  1.4041e-01,
         -6.2742e-02, -5.7964e-02, -1.7902e-01, -4.5360e-02, -8.5336e-02,
         -3.2277e-01, -3.3387e-01, -1.9794e-01, -1.0924e-01, -7.9379e-02,
         -1.7139e-01, -2.1645e-01,  2.8733e-02, -2.0589e-01, -1.3113e-01,
         -1.3366e-01,  3.9030e-02, -1.3969e-02,  5.3785e-02, -7.2571e-02,
          9.6827e-02,  5.6421e-02, -5.5339e-02,  2.7051e-02, -7.0325e-02,
          4.8131e-02,  8.1803e-02,  3.3510e-02,  1.7082e-01,  1.4118e-02,
         -5.3776e-02, -1.1917e-01, -1.3166e-01,  1.3488e-01,  3.8569e-02,
          2.0678e-01,  6.3014e-02, -1.6616e-01, -7.6079e-02, -9.8365e-02,
          1.0504e-01,  1.8116e-01,  1.0582e-01, -1.4959e-01, -8.6256e-02,
         -2.5763e-02, -1.5695e-02, -2.6077e-02,  4.7794e-02, -2.1334e-01,
         -7.0313e-02,  7.9473e-03,  1.3277e-02, -1.6328e-01, -7.7013e-02,
         -2.5627e-02,  9.2429e-02,  1.0088e-01, -2.7362e-03,  4.1562e-01,
          6.1893e-03,  1.4407e-01,  2.9154e-02,  1.2896e-01,  1.5596e-01,
         -9.8563e-02,  2.2995e-01, -2.8181e-02, -7.6099e-02, -6.3219e-02,
         -1.4815e-01, -1.9633e-03, -9.9625e-03,  2.0166e-01,  4.6836e-02,
          5.2547e-02,  1.8354e-01, -4.1396e-02,  1.6370e-01,  2.3645e-02,
          1.2548e-01,  8.2798e-02, -7.4780e-02,  1.2656e-01,  1.7083e-01,
          7.2788e-03,  6.7456e-02,  1.4332e-01, -4.4247e-02,  1.1582e-01,
         -1.7354e-01,  1.4678e-01, -4.8418e-02,  6.1749e-02, -1.1245e-01,
          1.6182e-03, -4.4248e-02,  2.1827e-02, -3.4436e-02,  2.2592e-02,
         -1.3858e-01, -1.3659e-01,  1.2117e-01, -4.2950e-02, -9.0023e-02,
         -1.2190e-02, -9.7948e-02,  2.9256e-02, -4.7738e-02, -1.1670e-02,
         -7.6813e-02,  8.5547e-02, -2.4177e-02,  1.1507e-02,  4.3484e-02,
         -1.0297e-01,  2.6449e-03,  1.3819e-02, -4.7608e-02,  2.0875e-02,
         -3.7713e-02, -1.2329e-01,  1.6512e-02,  1.5769e-01, -1.1697e-02,
          2.3357e-02,  5.2645e-02,  1.2846e-01, -6.7302e-02,  1.4715e-01,
          1.7625e-01, -3.2995e-02, -2.6747e-02, -5.5318e-02,  1.6758e-01,
          1.0104e-01,  1.1779e-01, -4.9764e-02, -8.2016e-02, -6.9898e-02,
         -5.9184e-02,  3.9349e-02,  3.8230e-03, -1.2207e-01, -4.4911e-02,
         -2.1776e-01, -1.5588e-01,  1.1355e-01,  1.6922e-01, -1.3374e-01,
          1.2142e-01,  3.4891e-03,  2.0870e-02,  7.4153e-02,  4.4189e-02,
          1.7416e-01, -7.3337e-02,  1.2243e-01, -1.1373e-01,  1.4150e-01,
         -7.6444e-02, -4.5403e-02, -1.1519e-01,  4.3861e-02,  6.6192e-02,
          3.2538e-02,  1.1703e-01, -1.2036e-01, -8.7026e-02, -7.0192e-02},
        '{-3.3784e-02, -9.9313e-02, -4.3042e-02, -8.6584e-02,  1.5053e-02,
          1.1633e-01,  1.1557e-01,  2.1181e-02,  1.0230e-01,  6.1452e-02,
         -3.2138e-02,  1.1588e-01, -4.3730e-02, -5.3300e-02, -1.2003e-01,
         -3.2171e-02, -2.0368e-02,  5.7392e-02, -1.1906e-01, -3.4288e-02,
         -1.9395e-02, -7.3425e-02, -1.1422e-01, -7.2927e-02,  3.3491e-02,
         -5.9271e-02,  7.3901e-02,  6.2827e-03,  1.9239e-02, -8.7586e-02,
          3.6394e-03, -2.0372e-03, -9.7463e-05,  1.8456e-02,  1.6124e-02,
         -2.1970e-03,  3.0126e-02,  6.7441e-03, -1.0052e-01,  6.8160e-02,
          3.5893e-02,  3.5226e-02, -3.6268e-02,  4.5245e-03, -5.3512e-03,
          9.4557e-02,  5.0290e-02, -4.9764e-02,  1.2208e-04, -5.0186e-04,
          4.2296e-03,  2.2728e-02,  1.9166e-02,  6.0148e-02,  3.2368e-02,
         -8.1354e-02,  3.7620e-03,  3.2422e-02, -4.3975e-02, -4.6835e-03,
         -4.7811e-02, -6.5291e-03, -1.0848e-01,  2.3108e-02, -3.8712e-02,
          1.1245e-01, -2.3701e-02,  1.9196e-02,  3.4154e-02, -8.6216e-02,
         -8.4216e-02,  9.2208e-02, -1.0162e-01, -8.1175e-02, -1.0873e-02,
         -5.0361e-04, -3.3394e-02, -4.5211e-03,  5.6951e-02, -2.1446e-02,
          1.9426e-03, -1.2324e-02, -1.1346e-02,  8.4866e-03, -6.3270e-04,
          7.4310e-03, -2.3970e-22, -4.3573e-03,  5.6979e-03,  1.5397e-02,
          2.9161e-03,  9.3138e-09,  3.1169e-03,  6.0485e-02, -2.4782e-02,
         -6.1714e-02,  8.6769e-03,  3.0093e-02, -5.1780e-02, -4.4953e-03,
          2.2538e-02,  7.7652e-02, -5.3051e-02,  7.4356e-02, -5.0948e-02,
         -2.5484e-03,  4.5769e-02,  8.2888e-02, -1.4893e-01,  6.8391e-02,
          1.9456e-02, -1.9268e-02,  5.2551e-02, -4.1148e-02, -1.7705e-02,
         -6.2490e-02, -1.3380e-01, -2.7558e-02,  1.2639e-03,  2.4973e-02,
         -1.5086e-02, -7.5776e-02, -5.7860e-03, -1.1876e-01,  1.0081e-01,
          3.2619e-02,  2.2719e-02, -7.1717e-03, -5.6424e-03, -3.8468e-02,
          2.0879e-06, -3.1764e-02,  5.5351e-02, -6.0693e-02,  3.3505e-02,
          3.6561e-02,  1.0093e-01,  4.4126e-02,  1.1506e-02, -8.2574e-02,
          4.0010e-02, -3.4217e-03, -1.3302e-02,  2.6268e-02, -2.9743e-02,
          3.3406e-02,  3.3679e-02, -7.2260e-02,  6.4361e-03, -3.5779e-02,
          1.4863e-02, -5.3570e-02,  1.0606e-02,  7.9166e-03, -6.4952e-03,
         -6.7991e-02, -1.5033e-01, -1.7534e-02, -9.9559e-02, -3.5710e-04,
          7.0737e-02,  9.3831e-02, -8.3267e-02, -3.4946e-02, -4.3209e-02,
          4.9801e-02,  5.7669e-02,  3.9606e-02,  5.4196e-03, -8.8438e-02,
          6.7013e-02, -9.9125e-04,  4.0199e-02, -3.3584e-02,  8.1938e-02,
         -6.1506e-02, -6.4570e-02, -2.3703e-02, -8.8414e-02,  2.6063e-03,
          1.1975e-01, -4.6478e-02,  1.2868e-01, -9.0698e-02, -9.0623e-03,
          5.3059e-02, -8.3291e-02,  2.5883e-02, -6.1827e-02, -1.1212e-01,
         -7.1555e-03, -2.2602e-02, -8.3120e-02, -5.6628e-02,  4.8283e-03,
         -8.5341e-02,  8.8716e-02, -9.8658e-02,  5.5309e-02, -1.1657e-03},
        '{ 3.8888e-03, -1.4028e-01, -1.2678e-03,  1.1009e-01,  4.9753e-02,
         -5.0538e-03, -2.7698e-02,  4.1762e-03, -1.1443e-01, -1.8970e-02,
          6.3849e-02, -6.1451e-02, -1.5938e-01, -2.4815e-01, -1.2879e-01,
         -6.8029e-02, -7.1407e-04, -3.6109e-02, -7.5408e-02, -1.9420e-02,
          2.3907e-01,  1.5180e-01,  4.9701e-02,  6.2702e-02,  1.2928e-01,
          4.6110e-02,  2.5389e-01,  1.5318e-01, -9.2358e-02, -7.7216e-02,
          8.0716e-02,  1.5186e-01,  1.0255e-02, -2.2326e-01, -1.3425e-01,
          1.8084e-01,  9.4949e-02,  6.3971e-02,  7.2861e-02, -1.9603e-02,
         -4.2096e-02,  5.7522e-02,  1.4444e-01, -3.8838e-02,  4.4974e-02,
         -1.4825e-02, -7.4491e-02,  1.1073e-01,  1.8034e-01,  6.8063e-02,
         -2.3587e-03, -1.1437e-01,  2.3787e-01,  2.4788e-02,  2.4153e-02,
         -9.7427e-02,  1.0622e-02,  1.5367e-01,  7.2994e-02, -2.9647e-02,
         -3.3743e-02, -2.7437e-02, -2.8345e-03,  8.2230e-03, -1.0466e-01,
          4.0090e-02, -8.2096e-02, -6.3956e-02, -2.2903e-01, -3.1597e-02,
          1.0464e-01, -1.4527e-01,  1.2375e-01,  1.1027e-01,  7.1869e-02,
          8.7502e-02, -3.4926e-02, -6.7300e-02, -3.5278e-02,  2.5637e-02,
         -2.7321e-02, -3.4597e-02,  1.0827e-01,  7.6559e-02,  6.8934e-02,
         -5.3330e-02, -9.5715e-02, -1.2382e-03,  6.6485e-02,  1.1956e-01,
         -3.9267e-03, -6.1153e-02, -7.7660e-02,  7.2278e-03,  8.7978e-02,
         -6.6139e-02, -3.3093e-02,  1.9103e-02,  6.5084e-02,  2.2314e-02,
          4.1630e-02,  1.2488e-02, -1.0420e-01,  1.9374e-01,  9.9322e-03,
         -9.3938e-02, -1.0950e-01,  1.0873e-01,  1.5261e-01, -7.7131e-03,
          1.5272e-01, -1.1393e-01, -3.1799e-02, -1.0340e-02, -1.8079e-01,
         -1.0126e-02, -6.2278e-02,  8.0312e-02,  5.4898e-02,  1.1562e-01,
          1.7200e-01,  7.5774e-02,  1.2858e-01, -1.1108e-02,  1.2723e-01,
          4.9870e-02,  2.2115e-01,  3.7847e-02, -1.6168e-01, -3.5556e-02,
          1.8444e-01,  1.3417e-01,  9.6087e-02, -9.0953e-02, -1.7045e-01,
          8.4484e-02, -1.2201e-02, -8.0026e-02,  3.9957e-02, -2.9502e-02,
         -8.7638e-02, -1.1002e-01, -1.2060e-01, -1.3292e-01, -9.0349e-02,
          6.7860e-02,  1.3368e-01, -6.3111e-02,  2.1272e-01,  1.6283e-01,
         -3.3349e-02, -4.0509e-02, -5.1881e-02,  7.8040e-04, -4.0426e-02,
          3.7104e-02,  7.3259e-02, -3.6849e-02, -1.0962e-01,  9.3134e-02,
         -6.6259e-02,  3.4450e-02,  9.0986e-02, -1.8013e-01, -6.6425e-02,
          7.5730e-02, -1.1195e-01,  1.2875e-01, -4.9576e-03,  1.1036e-02,
          8.9207e-02, -8.6124e-02,  5.6901e-02,  1.0285e-01,  7.3701e-02,
         -9.4986e-02,  1.2968e-01, -1.1773e-01,  2.0656e-02, -3.9925e-02,
         -1.0561e-01,  5.1201e-02,  4.1048e-02,  1.5975e-01, -7.5954e-02,
          8.1237e-02, -1.2163e-01,  4.2089e-02, -1.4281e-01, -6.0320e-02,
          1.1034e-01,  1.5172e-01,  8.9191e-02, -1.5078e-02,  2.5815e-02,
         -5.2166e-02,  1.2571e-02, -4.4428e-02,  1.1394e-01,  1.9449e-01},
        '{ 1.7129e-01, -1.2413e-01, -8.6345e-02, -1.3191e-01,  8.6816e-02,
         -5.2373e-02, -1.2758e-01, -1.7362e-01,  3.1744e-03, -1.4710e-01,
          6.6178e-02,  9.3161e-02,  1.3795e-01,  5.4334e-02, -1.3807e-01,
         -1.1922e-01,  1.0323e-02,  8.0247e-02,  7.8893e-02,  1.7169e-01,
         -2.0585e-01, -1.9764e-01, -1.0976e-01,  1.7912e-01,  2.5129e-02,
         -1.1155e-02, -3.0472e-02, -6.7915e-02, -1.9806e-01, -1.1018e-01,
          1.5605e-01, -6.5269e-02, -1.5439e-01, -3.3464e-01, -8.2578e-02,
          6.2537e-02,  7.7258e-02, -6.6863e-02, -1.6187e-01,  1.0983e-01,
          3.7922e-02, -3.3189e-02,  1.8979e-02, -7.4697e-02, -1.1183e-02,
         -1.4331e-01, -1.0234e-01, -3.9510e-02, -6.6779e-02,  1.8114e-01,
          7.6725e-02,  5.1070e-02,  5.5221e-02,  1.6188e-01,  1.7625e-01,
          3.1673e-02,  1.0185e-01, -8.6798e-02, -1.2342e-01, -6.2577e-02,
          6.9403e-02,  1.9662e-02,  7.4306e-03, -3.4855e-02, -1.1258e-01,
          1.1134e-01,  6.7946e-02,  3.4242e-02,  3.7141e-02, -3.3976e-02,
          4.7468e-02,  8.2791e-02, -7.0135e-02,  6.1106e-02, -4.0679e-02,
         -2.8278e-02, -2.9721e-02,  1.0553e-01,  2.6083e-01,  8.4977e-02,
         -1.0722e-01, -8.4707e-02,  7.1986e-02,  1.9514e-01,  3.3275e-01,
         -8.6555e-03,  8.0839e-02, -6.3932e-02, -8.9227e-03,  1.1356e-01,
          1.8473e-02,  1.5658e-01,  2.1867e-01, -1.8593e-02, -1.0369e-01,
          1.2090e-01,  1.4418e-01, -1.1925e-01,  1.4688e-02, -1.6049e-01,
          8.5117e-02,  7.3472e-02,  1.5237e-01, -3.9504e-02,  1.1797e-01,
         -1.1314e-01, -7.6333e-02, -2.8131e-04,  6.0657e-02, -1.2609e-01,
         -1.1014e-02, -1.0524e-01,  1.5563e-01,  8.6745e-02,  3.7320e-02,
         -1.1313e-01,  8.0469e-02,  3.2230e-02,  6.7123e-03,  5.9624e-02,
          4.8307e-02,  8.3660e-02, -5.2053e-02, -9.3103e-02,  8.9850e-02,
         -9.3340e-02,  1.1054e-01,  1.8237e-01, -4.8191e-03,  7.9853e-02,
          1.2400e-01,  8.5544e-02, -8.1937e-02, -2.3499e-01, -1.8044e-01,
         -1.3114e-02,  9.1901e-02,  4.4341e-02,  5.9347e-02, -4.9330e-02,
         -3.1058e-02, -3.8668e-02,  1.3256e-01,  1.6092e-01, -2.7658e-02,
         -1.9416e-02,  1.4291e-01,  1.7440e-02,  1.1313e-01, -8.3919e-02,
         -4.8845e-02,  1.3004e-01,  1.3580e-01, -4.9343e-02,  1.0617e-01,
         -5.1377e-02,  7.9908e-02, -7.8227e-02,  6.9238e-02,  1.5938e-01,
          1.1044e-01,  1.9723e-03,  1.6626e-01,  1.3193e-01, -4.5978e-03,
          1.2340e-01,  2.1620e-03,  1.6958e-01, -1.6412e-02, -7.0438e-02,
          9.3788e-02, -1.0703e-01, -1.1726e-01, -1.1685e-01,  5.3299e-02,
          1.1910e-01,  4.9561e-02, -9.5053e-02, -1.9833e-02,  2.9120e-02,
          1.2126e-01, -7.0024e-02,  1.1679e-01,  1.2975e-01, -1.2000e-01,
         -8.9582e-02,  6.1831e-02,  6.7533e-02, -7.4769e-02, -2.3765e-02,
          1.1114e-01,  1.3842e-01,  1.8088e-01,  5.0120e-02,  6.6975e-02,
          8.4727e-02, -1.0299e-01,  1.0324e-01,  7.1807e-02, -7.3689e-02},
        '{-1.3368e-01,  4.2059e-02,  6.8800e-02, -6.6091e-02, -8.7037e-02,
         -6.2383e-02, -7.8442e-02,  1.4772e-02,  1.3285e-02, -5.3030e-02,
          8.1768e-02,  2.4030e-02, -2.2771e-01, -2.1462e-01,  4.7626e-02,
          1.0883e-02,  9.3946e-02, -1.1730e-02,  1.0655e-02, -9.9579e-02,
         -1.3465e-02, -3.0138e-02, -9.1989e-03, -1.0205e-01,  4.3332e-02,
         -8.9641e-02,  3.5074e-02, -4.0884e-02, -5.9869e-02, -3.1019e-02,
          5.9966e-02,  3.3012e-02, -2.3139e-02,  8.0902e-02,  8.3138e-03,
         -8.1502e-02, -1.1609e-01,  5.1597e-02,  1.3891e-01, -2.4565e-01,
         -1.6452e-01,  2.9463e-03, -4.8267e-02,  9.5215e-02, -6.5051e-02,
         -4.1686e-02,  8.3816e-02,  1.1141e-01, -2.3476e-02,  1.7058e-01,
          1.1824e-01,  4.4456e-02, -7.9564e-02,  1.0751e-02,  6.3107e-02,
          1.2075e-01, -3.5941e-03,  2.0816e-02, -8.6926e-02,  9.6761e-02,
          4.3506e-02,  6.3758e-02, -1.0733e-01,  1.4556e-01,  1.7326e-01,
          1.4768e-01, -2.4111e-03,  4.2348e-03, -1.0073e-01,  9.3797e-02,
         -8.5820e-03,  1.2915e-01, -1.5425e-02, -1.1698e-01, -9.2105e-02,
          4.1358e-02, -5.7269e-02,  3.9418e-02,  5.7530e-02,  4.7447e-02,
         -7.8630e-02,  1.4136e-01,  1.3193e-01,  1.7814e-01, -4.0212e-02,
         -2.0025e-02, -1.0424e-01,  1.0579e-01,  1.3030e-01,  7.3078e-02,
         -1.0065e-01,  1.9045e-01,  6.3112e-02,  5.4131e-02,  1.2416e-01,
          7.3581e-02,  1.2442e-01, -1.7684e-02,  1.1082e-02, -1.6178e-01,
         -1.0500e-01,  1.1868e-01,  2.2844e-02,  1.4174e-01, -7.9621e-02,
          1.3637e-01, -3.5488e-02,  9.5018e-02,  1.1559e-01, -3.2922e-02,
          7.4184e-02, -3.3059e-03, -6.5362e-02,  3.4206e-02,  2.7870e-02,
         -8.6390e-02,  1.4365e-01,  9.1406e-02,  1.2446e-01,  2.0220e-02,
         -6.2832e-02,  1.8883e-01,  1.3514e-01, -1.9433e-02,  1.8449e-01,
          3.9391e-04, -4.2070e-02,  7.0963e-02, -2.4573e-02,  1.1510e-01,
         -2.1781e-03, -1.3900e-02,  1.1002e-01,  1.6231e-01, -5.5813e-02,
         -1.1381e-01, -1.9357e-01, -1.0009e-01,  3.2148e-03, -2.6656e-02,
          8.9525e-02, -1.7034e-01, -1.5292e-01, -1.6191e-01,  1.6624e-01,
          2.0002e-02, -8.7042e-02,  1.1989e-02,  1.1801e-01,  5.3937e-02,
         -1.2016e-02, -1.4233e-01,  2.2147e-02,  6.6603e-02, -1.1070e-01,
          8.4789e-03,  4.1036e-03,  1.3033e-01, -1.2292e-01, -5.8714e-03,
          1.3807e-02,  8.2450e-02, -1.7289e-01, -9.8865e-02,  3.7045e-02,
          3.7512e-02,  8.9899e-02,  7.4673e-02,  1.5593e-01,  7.9276e-02,
         -1.0764e-01,  1.4461e-01,  1.8253e-01, -1.1583e-01, -9.2449e-02,
         -1.0239e-01, -5.7501e-02, -1.2269e-01, -9.5771e-02, -1.5278e-01,
         -1.4523e-02,  1.1002e-01, -1.1489e-01,  1.3916e-01,  2.2533e-02,
          1.0580e-01,  8.0267e-02, -1.6692e-01, -1.5628e-01,  1.6636e-01,
          1.4395e-01,  2.1368e-01,  1.1474e-01, -1.7773e-02,  1.1042e-01,
         -1.5550e-01, -9.2433e-02,  1.7543e-01, -1.0945e-01, -4.2176e-02},
        '{-1.0139e-01, -1.5144e-01,  1.1525e-01, -3.2459e-02,  9.1015e-02,
         -9.8071e-02, -1.9189e-02,  6.1899e-03,  1.5670e-01,  1.1985e-01,
         -9.2654e-03,  8.9871e-02,  2.0769e-01,  1.5271e-01,  1.0146e-01,
         -3.9065e-02, -2.4182e-02, -5.7055e-02,  4.6717e-02, -1.7003e-01,
          7.3936e-03,  1.3758e-01,  4.2875e-02,  9.5612e-02, -1.4870e-01,
         -7.2297e-02,  1.0938e-01, -2.2717e-01,  2.6937e-02,  3.5164e-02,
         -5.8109e-02, -3.8563e-01, -1.5588e-01, -1.0381e-01,  2.4816e-01,
         -1.3623e-01, -3.7250e-02, -6.9692e-02,  1.2472e-01,  1.3687e-01,
         -4.1301e-02, -9.2988e-03,  1.7305e-01, -5.5520e-05, -5.8075e-02,
          4.5651e-02,  8.4591e-02, -8.1239e-02, -6.7539e-02, -4.0766e-02,
         -1.2006e-01,  9.8116e-02, -7.4894e-02, -1.0384e-01, -2.5185e-01,
          2.5882e-02, -1.2569e-01,  6.9765e-02,  8.6216e-02,  1.5685e-01,
          1.1244e-01,  2.0110e-01,  9.1643e-02,  1.5616e-02,  2.0109e-01,
         -1.3568e-01, -3.4713e-02,  5.9237e-02,  2.6881e-02,  1.4577e-02,
         -1.8625e-02, -5.6125e-02, -8.5159e-03, -2.1386e-03, -2.0608e-01,
         -1.7539e-01, -7.6634e-02,  1.1785e-01,  8.2333e-02, -2.9400e-02,
         -4.4879e-02, -8.0493e-02,  8.0758e-02, -2.1038e-01, -8.9179e-02,
         -1.0979e-01,  1.1596e-01, -4.4570e-02, -2.4584e-01, -8.4768e-02,
         -1.2090e-01, -3.0054e-02, -5.7731e-02, -1.1997e-01, -6.3986e-02,
          7.2544e-02,  5.8765e-02,  7.8488e-02, -9.5680e-03,  6.2626e-02,
         -7.6362e-02,  7.2622e-03,  1.3660e-01, -8.6765e-03,  1.1974e-01,
         -1.6279e-01, -8.0094e-02,  1.6259e-01, -1.1857e-01, -1.1647e-01,
          3.1882e-02, -1.1456e-01, -2.2972e-02,  1.8619e-02, -1.4764e-01,
          6.1469e-02, -9.5257e-02,  8.7866e-03,  6.4963e-02, -5.0369e-02,
         -8.2085e-03,  8.4447e-02,  1.2699e-01,  1.5089e-01,  1.1335e-01,
         -9.8408e-02, -1.3973e-01, -2.3050e-01, -7.9706e-02,  2.2771e-01,
         -1.7549e-01, -6.0072e-02,  2.6136e-02, -3.6966e-03,  1.4193e-02,
          1.3471e-02,  7.0078e-02,  1.4979e-01, -3.7185e-03,  1.9312e-01,
         -1.1516e-01,  1.2407e-02,  2.3398e-03,  6.9443e-02, -2.1616e-01,
         -8.9941e-02,  1.0291e-01, -6.2432e-02, -1.2806e-01, -1.1794e-01,
          1.3815e-02,  6.2525e-02, -5.6779e-02, -1.3053e-02,  1.4191e-01,
          9.7837e-02, -8.2879e-02, -1.2495e-03, -4.1501e-02, -1.2125e-01,
         -1.6031e-01,  7.9664e-02,  4.7518e-02,  1.8006e-01, -1.3159e-02,
         -3.3746e-02, -1.4759e-01, -9.9764e-02,  3.3560e-02, -3.4197e-02,
         -1.5548e-01, -3.3036e-02,  1.5882e-01, -7.9778e-02,  9.2575e-03,
         -8.5513e-02, -1.5286e-01,  3.1384e-02,  7.7025e-02, -1.0528e-01,
         -1.4188e-01,  1.5483e-02, -2.6398e-02,  5.9787e-02, -1.3245e-02,
         -4.5697e-02, -1.1542e-01,  1.4981e-01, -7.3523e-02,  2.1625e-02,
         -4.6224e-03,  9.7181e-02, -1.5600e-02, -2.7093e-04, -2.0930e-01,
         -1.2658e-01,  8.3817e-02,  1.3576e-01,  7.4259e-02, -1.1791e-01},
        '{-9.3511e-02,  3.3892e-02, -1.7802e-03, -4.7684e-02,  7.5975e-02,
          7.8440e-02, -1.3124e-01, -8.8813e-02,  7.8802e-02,  1.4555e-01,
          2.5093e-02, -5.6102e-02,  7.5143e-02, -2.4821e-02,  1.7613e-01,
          1.4329e-01, -1.0198e-02,  1.5213e-01,  4.5266e-02,  1.2812e-01,
         -1.5657e-01, -5.9008e-02,  1.0123e-01, -5.2944e-02, -5.5187e-02,
          9.9764e-02, -3.2258e-02,  4.3386e-02,  4.4522e-02,  1.0260e-01,
         -7.9341e-02, -1.1251e-01,  5.0619e-02,  6.6253e-02,  7.3860e-02,
         -2.5016e-01, -2.1216e-01, -3.2471e-02,  1.7395e-01,  9.3774e-02,
          6.0294e-02, -1.1380e-01, -1.5974e-01,  8.2791e-02,  1.7416e-01,
         -5.2480e-02, -8.7337e-02,  2.7176e-02, -1.0100e-01, -5.4213e-02,
         -4.6104e-02,  6.9002e-02,  8.4588e-02, -1.8174e-02,  6.6444e-02,
         -9.8792e-02, -2.7721e-03, -1.4048e-01,  3.2014e-02, -9.8754e-02,
          6.9065e-02, -2.1378e-02,  5.4669e-02, -4.0660e-03,  2.5977e-02,
          1.3437e-01,  5.4203e-03,  4.6385e-02,  8.7049e-02,  4.8894e-02,
         -7.0230e-02,  8.6744e-02,  1.4071e-01, -1.1992e-01, -7.9797e-02,
          1.9708e-02,  2.2213e-02,  1.2704e-01,  4.7895e-02,  1.4551e-01,
         -1.0542e-01, -4.7683e-02,  5.0623e-02, -5.1479e-02,  3.9319e-02,
         -2.4645e-02,  1.1771e-01, -2.0272e-02, -1.1285e-01, -9.0443e-02,
         -2.7454e-02, -8.8556e-02, -7.2037e-02,  1.5959e-01, -1.2690e-01,
         -2.5910e-02, -8.7630e-02,  1.6104e-01,  3.9452e-02,  1.0697e-01,
          1.2040e-01, -3.5209e-02, -1.4818e-02,  3.8249e-02, -7.1432e-02,
         -1.4173e-02,  1.5494e-02,  8.8566e-03, -4.2325e-02,  3.0200e-02,
          8.8368e-02,  8.5349e-02, -1.5774e-01,  3.6971e-02,  1.4742e-01,
          5.7600e-02,  3.1087e-02, -7.4791e-02, -3.8035e-02,  2.8008e-02,
          3.9863e-02, -3.3175e-02, -1.2553e-01,  9.0414e-02,  4.7088e-02,
          7.5238e-02, -2.3072e-01, -7.3653e-03, -8.6430e-02, -1.2503e-02,
         -8.2378e-02, -1.1662e-01,  5.3345e-02,  7.6891e-03,  2.3113e-01,
         -1.2691e-01,  1.3349e-01, -3.4134e-02, -5.8040e-02, -2.2932e-02,
          3.8829e-02,  3.4272e-02, -4.3039e-02, -1.7010e-02,  1.3630e-01,
          2.5606e-02,  3.5022e-02,  4.7418e-02,  1.9611e-02,  4.8436e-02,
         -7.6803e-02, -2.8807e-03,  8.1354e-02,  4.9830e-02,  1.6543e-01,
         -4.3414e-02,  1.4492e-02,  1.3256e-01,  9.2643e-02, -9.4373e-03,
         -8.8553e-02, -1.2864e-02, -1.1302e-01, -9.4026e-03,  3.0529e-02,
          5.5819e-02,  8.6146e-02, -1.3455e-01,  6.1752e-03,  1.5531e-01,
         -8.2836e-02, -9.4333e-02, -1.5526e-02,  1.2568e-01,  4.5297e-02,
         -9.2038e-02,  1.2367e-01, -1.8395e-01,  5.6392e-02,  9.0614e-02,
          3.0719e-02,  2.0355e-01, -6.7645e-02, -9.5512e-02,  4.7863e-02,
          1.1446e-01, -2.7521e-02,  2.7607e-02,  3.9400e-02, -3.3112e-02,
         -3.6824e-02,  7.0326e-02, -2.4088e-02,  7.5208e-02,  1.1029e-03,
          1.0072e-02,  8.8814e-02,  1.9253e-02,  3.9317e-02, -8.3051e-02},
        '{ 1.5814e-01, -1.0721e-02, -1.0303e-01, -7.1254e-02,  1.8423e-02,
         -3.9852e-02, -8.2209e-02,  8.4128e-02,  1.0289e-02,  7.0049e-02,
          1.4304e-01,  2.5214e-02, -5.0801e-02,  1.2460e-01,  6.7076e-02,
          1.7279e-01, -8.9770e-03,  5.8061e-02,  1.5182e-01, -1.5421e-02,
          9.8658e-02, -1.8913e-01, -1.2207e-01, -7.3742e-02,  2.6373e-01,
          1.9748e-01,  9.7285e-02,  6.8986e-02,  1.8284e-01, -2.1814e-02,
          3.2711e-01,  1.0772e-01,  1.6285e-01,  6.2640e-02, -1.1461e-01,
          1.1183e-01,  1.6118e-01,  7.0740e-02, -1.0587e-01, -7.3608e-02,
          1.7043e-01, -6.1148e-02, -4.8975e-02, -4.8346e-03,  2.6105e-01,
         -4.5354e-02, -7.2738e-02,  1.0933e-01,  5.5170e-03,  1.8787e-01,
          1.1235e-02,  1.4045e-01,  3.4228e-02,  2.1161e-01,  1.2690e-01,
         -1.1035e-01,  7.6840e-02,  2.5640e-03, -1.0808e-01, -4.2882e-02,
         -6.2743e-02, -1.4326e-01,  1.3367e-01, -3.9793e-02,  3.8041e-02,
         -4.6906e-02, -9.5496e-02,  8.7115e-02, -6.4805e-02,  8.7579e-02,
         -1.2556e-01,  4.0550e-02, -5.2404e-02, -3.4591e-02,  2.7905e-02,
         -2.7958e-02, -5.8916e-02, -2.2090e-02,  5.0349e-02,  3.7416e-02,
         -1.0237e-01, -1.1305e-01, -4.1221e-02,  1.7513e-02,  4.8212e-04,
          8.0801e-02, -1.3531e-01,  9.8036e-02, -4.6022e-02, -1.4065e-02,
         -8.7651e-02,  1.1402e-01,  1.8296e-01,  6.6826e-03,  3.5752e-02,
          6.8520e-02,  4.4981e-02,  1.4896e-01, -4.4882e-02, -1.3565e-01,
         -6.1432e-02, -9.4001e-02, -6.8392e-02,  1.6812e-02, -3.6706e-02,
          1.1242e-01, -8.1175e-02, -1.0203e-01,  8.4462e-02, -1.7525e-01,
          1.9779e-02, -7.1569e-02,  6.1911e-02, -1.0202e-01,  1.3143e-01,
         -6.2694e-03, -2.4217e-03,  2.0651e-01,  9.9633e-02, -1.3176e-01,
          1.8069e-02,  1.7072e-01, -2.6276e-02,  9.2894e-02,  3.7932e-02,
          6.9141e-02,  2.4698e-02, -4.1436e-02,  1.5805e-01,  1.2689e-01,
          1.6130e-01,  1.0725e-01,  2.0427e-01, -1.1522e-01, -3.0118e-02,
          4.2213e-02,  6.2459e-02, -1.2670e-01,  6.3470e-02, -7.8973e-02,
          1.0777e-02,  9.1544e-02,  3.5427e-02,  8.6868e-02,  1.2718e-01,
         -6.4976e-03,  6.8605e-02, -7.7692e-02, -3.1694e-03,  8.0318e-02,
         -3.2481e-02,  1.4791e-01,  1.4051e-01, -1.3452e-01, -1.4685e-01,
          1.5011e-01, -1.0306e-01, -5.6862e-02,  1.5582e-01,  3.3147e-02,
         -1.1722e-01,  1.1634e-01,  9.0882e-02,  1.8466e-01,  1.0262e-01,
         -1.2531e-02,  1.0481e-01,  1.9376e-02,  1.2332e-01,  3.3110e-02,
          1.4410e-01, -3.0832e-02, -5.9356e-02, -9.6623e-02,  8.8556e-02,
          1.1253e-01,  3.4985e-02, -2.1069e-02,  5.1797e-02, -4.5710e-02,
          6.2899e-02, -1.5852e-01,  2.1990e-02,  1.5046e-02,  5.7911e-02,
         -1.2581e-01, -2.6650e-02,  6.3346e-02,  2.2011e-02, -5.0715e-02,
          1.3790e-01,  4.4815e-02,  1.3400e-01,  7.2357e-02,  8.8723e-02,
         -9.1415e-02, -8.3517e-02,  9.3702e-02,  1.1868e-01,  1.3410e-01},
        '{-1.0397e-01,  3.0090e-02,  1.0168e-01,  1.0226e-01,  1.6303e-02,
          7.8107e-02, -1.1319e-01, -7.7299e-03, -2.1850e-03, -4.3292e-02,
         -1.2248e-01,  5.8393e-02,  6.4606e-02,  1.2778e-01,  6.7951e-02,
          8.5541e-02,  1.5635e-01,  2.0818e-02,  1.0590e-01, -5.6840e-02,
          1.4486e-02,  6.0613e-02,  1.0967e-01, -2.2604e-02,  3.0676e-02,
         -4.3899e-02, -8.3204e-02, -1.0219e-01, -1.2637e-01, -1.2808e-01,
         -1.0356e-01,  1.4896e-02, -1.0188e-01, -2.1492e-01,  9.7098e-02,
          1.3594e-01, -1.4347e-02, -1.2078e-01,  1.9463e-01, -5.8393e-04,
         -7.9796e-02, -4.6007e-02,  2.3089e-02,  6.8216e-02, -1.3894e-01,
         -3.5143e-02, -2.6755e-02,  1.0173e-01,  1.1288e-01,  9.3115e-02,
         -1.0359e-01, -7.4307e-03,  9.6999e-02,  6.3616e-02, -3.9957e-02,
         -7.4015e-02, -8.2372e-03,  1.1411e-01, -6.7120e-02,  5.5472e-02,
          3.8692e-03, -3.5934e-02,  4.4747e-02, -6.4488e-02,  1.3868e-02,
         -1.4778e-01,  2.0056e-02, -7.1544e-02,  1.5727e-01, -3.9527e-02,
         -1.4040e-02,  9.3189e-02,  1.0136e-01, -5.9240e-02, -1.2425e-01,
          1.5685e-02,  8.5562e-03, -1.9865e-02,  9.1865e-02,  5.5229e-02,
         -2.8906e-02,  7.1577e-02, -1.3098e-01,  1.6168e-01, -9.1557e-02,
         -1.9588e-02, -5.6741e-02,  5.4768e-02, -8.3469e-02, -2.5343e-01,
          3.0889e-02, -1.3536e-01,  1.3999e-01, -1.0979e-01, -7.7516e-02,
          5.9714e-02, -1.1129e-01, -7.8672e-02,  2.8993e-03, -2.0219e-02,
          1.4903e-01,  9.6423e-02,  1.0644e-01,  3.4784e-03,  1.3230e-01,
         -2.7791e-02,  2.9450e-02, -1.8155e-02, -9.8303e-03, -4.0899e-02,
         -1.3301e-02,  3.1000e-02, -3.8438e-02, -9.4112e-02, -1.8396e-03,
         -2.0913e-02,  4.1775e-02,  2.5120e-02, -1.2581e-01,  5.4730e-02,
          7.5804e-05, -5.3883e-02, -1.2516e-02, -3.1624e-02, -1.2434e-01,
         -7.9015e-02, -5.0014e-02,  1.3023e-01,  1.7939e-01,  8.9526e-02,
         -6.2494e-02,  4.8042e-03, -1.7271e-01,  6.9447e-02,  7.4360e-02,
          2.4842e-02,  2.7276e-02,  1.6916e-01,  1.6296e-01,  2.1239e-01,
         -7.4904e-02,  6.5163e-03,  1.0122e-01,  8.1317e-02, -5.7958e-02,
         -2.9021e-02,  4.5993e-02,  5.9628e-02,  9.7763e-03, -4.1594e-02,
         -9.7032e-02,  8.1986e-02,  1.2423e-02,  1.3318e-01, -1.2076e-01,
         -3.9720e-02,  9.0058e-03, -2.8448e-02, -1.5738e-02, -3.2114e-02,
         -7.3113e-03, -1.4247e-01,  1.4439e-01, -3.3737e-02, -6.3148e-02,
          5.8404e-02,  1.9680e-02, -2.5630e-02,  3.4683e-02, -4.0448e-02,
          1.3842e-01, -1.5542e-01, -4.1481e-02,  1.1759e-01,  2.8889e-03,
          9.6789e-02,  2.3862e-02, -1.5912e-02, -6.1803e-02, -2.6516e-02,
         -3.8920e-02,  6.5761e-02, -1.0999e-01,  1.1857e-01,  8.4824e-02,
         -3.9656e-02,  8.0862e-02, -9.5124e-02, -3.0468e-02, -1.5020e-01,
         -1.8007e-02, -9.3433e-02,  6.8159e-02,  9.5916e-02,  4.0219e-02,
         -8.9436e-03, -2.5803e-02, -1.6309e-01, -2.7586e-02, -3.5424e-02},
        '{ 3.3591e-02, -3.2983e-02,  3.2816e-02,  1.2084e-01, -8.2644e-02,
          9.6269e-04,  1.0004e-01, -8.2023e-02, -4.6509e-02,  9.4186e-02,
         -5.2490e-02, -1.5202e-02,  4.1241e-02, -6.1650e-02,  1.5422e-02,
         -2.3259e-02,  3.0171e-03, -1.2802e-02, -9.8124e-02, -8.1348e-02,
         -8.2149e-02,  1.1306e-01,  5.1870e-02, -1.4264e-02, -4.5247e-02,
         -1.5064e-01, -8.7215e-02, -1.0944e-01, -6.6003e-02, -9.3535e-02,
         -2.5259e-01, -3.7779e-03,  6.6551e-03, -1.3289e-01, -8.4149e-02,
         -3.2235e-01, -1.5579e-01, -2.0752e-01,  1.1226e-01, -2.3878e-01,
         -1.5704e-01, -3.3200e-01, -1.9234e-01, -2.1049e-01, -1.8340e-01,
         -1.4922e-01,  1.4420e-01,  6.7391e-02,  5.6131e-02,  9.7685e-02,
         -1.1250e-01, -3.6262e-02, -6.9459e-02,  8.4700e-02,  5.2326e-02,
          1.1455e-01, -3.8414e-02, -1.4902e-01,  3.6766e-03,  4.4927e-02,
          1.7149e-01, -8.4519e-02, -2.6834e-02, -1.8309e-02,  1.0641e-01,
         -3.5403e-02, -5.5725e-02, -8.3758e-02,  2.6137e-03,  7.9066e-02,
          1.3360e-01,  1.2726e-01,  1.3984e-01, -1.8143e-01, -1.3150e-01,
         -5.3995e-02, -5.6027e-02, -4.5099e-02, -1.5528e-02,  8.2294e-03,
         -8.9777e-02, -1.0322e-01, -3.6005e-02,  1.5340e-01,  2.2006e-02,
         -5.3224e-02,  1.3065e-01,  1.1863e-01,  7.3081e-02,  2.1577e-01,
         -6.9344e-02,  1.6196e-01, -6.2485e-02,  1.7259e-01,  1.8933e-01,
         -7.4759e-02,  1.8032e-02, -9.5460e-02, -1.4707e-01, -1.1170e-01,
         -8.3752e-03, -1.4118e-01, -1.1447e-01,  7.2054e-02, -1.9319e-02,
          1.2151e-01, -5.7145e-02,  1.3654e-01, -1.2217e-01,  1.6950e-02,
         -3.2169e-02,  1.3963e-01,  1.1905e-02, -1.1130e-01,  1.9349e-01,
          3.0320e-02, -7.6457e-02, -1.1620e-01, -2.8614e-02,  1.8394e-01,
         -1.1695e-01,  1.3131e-01,  1.0992e-01,  1.4120e-01, -1.4530e-01,
         -2.9889e-02, -1.3743e-02, -6.0539e-02, -1.2062e-01, -1.0372e-01,
         -1.1259e-01, -1.2607e-01,  4.4178e-02,  5.8324e-02, -6.0764e-02,
         -8.3110e-03, -1.3630e-01, -1.2257e-01,  1.1117e-01, -9.8406e-02,
          2.2320e-03, -1.5242e-01, -3.2014e-02, -6.7874e-02,  1.1199e-01,
          4.2204e-02,  1.1754e-01,  1.1455e-01, -7.9596e-02, -5.7010e-02,
         -1.3045e-03, -9.1763e-02,  1.1262e-01, -1.6740e-02, -9.3150e-02,
          4.4749e-02,  1.3370e-01, -4.3816e-02,  1.0403e-01,  1.2505e-01,
         -5.4035e-02,  1.4375e-01, -1.3839e-01, -5.4798e-02, -5.5806e-03,
         -3.4825e-02, -7.6116e-02, -1.2593e-01,  6.2977e-02,  1.5856e-01,
         -6.0857e-02,  3.1197e-02,  1.4099e-01,  1.6835e-01, -8.2823e-02,
         -1.1540e-01, -4.8780e-02,  7.7906e-02,  1.2716e-01, -1.7141e-02,
          5.3854e-02, -1.3586e-01,  1.9117e-02, -1.2486e-01, -5.4187e-02,
          2.1067e-01,  3.8926e-02,  5.5433e-02,  3.9525e-04,  1.0900e-01,
         -7.6867e-02,  1.4616e-01,  2.7147e-02,  8.7227e-03,  2.7064e-02,
         -2.1348e-02, -1.1341e-01,  3.0185e-02,  3.5845e-02,  5.4378e-02},
        '{-7.1825e-04,  1.3850e-02, -2.8838e-02, -5.2483e-02,  3.7426e-02,
          6.3718e-03, -5.1689e-04,  1.8610e-02, -3.0139e-02,  5.7537e-02,
         -1.2822e-02,  1.2003e-03,  7.7797e-02,  1.3020e-02,  6.4623e-05,
          2.6244e-02, -1.6037e-02, -2.2332e-02, -1.9618e-02,  1.7198e-02,
          6.6222e-02,  2.8434e-02,  1.0296e-02,  1.7152e-02, -7.0102e-03,
         -5.9220e-03, -1.4224e-02, -9.4672e-04, -1.5467e-02,  2.6882e-08,
         -6.4354e-04, -6.0398e-03, -2.2985e-05,  7.0627e-03, -4.4838e-02,
         -5.3987e-03,  1.1138e-09,  3.3946e-02, -1.4384e-02,  2.2658e-02,
         -2.5173e-05, -5.2463e-03,  1.7005e-02, -1.2114e-02, -3.7338e-03,
          2.6188e-03, -8.6059e-03,  3.8138e-08, -1.5513e-03, -3.3918e-02,
          1.9488e-03,  7.0457e-03, -1.5070e-03,  3.8293e-03,  1.4904e-02,
         -2.6554e-04, -2.4490e-02, -7.6093e-04,  2.7543e-02, -1.0538e-02,
         -8.5870e-03, -1.4943e-03, -9.6376e-04, -3.4358e-02, -2.8919e-02,
         -4.7008e-02, -1.5806e-03, -1.0339e-03, -9.4525e-03, -4.9222e-03,
          2.7134e-02, -5.1401e-02, -1.1801e-02,  1.5831e-02, -1.0953e-03,
          1.8830e-04,  2.3606e-02,  4.8648e-02, -3.6634e-02, -1.3331e-02,
          8.6469e-05, -7.0852e-03,  4.8338e-02,  2.5889e-03,  9.8529e-04,
          1.1859e-03, -5.2924e-02, -1.3365e-03,  3.5427e-03, -2.8547e-11,
          4.1930e-02, -1.5699e-03, -7.4247e-08,  3.1885e-03,  5.2426e-03,
         -3.8715e-02, -3.8203e-02,  1.8010e-03,  2.9655e-02, -7.1822e-04,
          2.2864e-03,  2.2001e-02,  4.8218e-02,  3.1786e-02, -3.4309e-03,
          3.5834e-03, -4.5041e-02,  3.5556e-02, -1.1055e-02,  6.4350e-02,
         -4.2295e-02, -1.0343e-03,  4.4987e-03,  4.2142e-02, -4.4324e-02,
         -6.5386e-02, -5.8194e-03, -2.2302e-02,  1.1198e-02, -9.9542e-03,
         -2.8596e-02, -7.6754e-02, -2.1282e-02, -1.7863e-03,  7.6844e-02,
         -5.2120e-04,  2.8149e-03, -2.0037e-03,  4.8213e-02, -1.6190e-03,
          6.6994e-04,  9.4291e-03, -2.5157e-02, -5.2853e-03, -7.0057e-02,
          4.7936e-05, -2.2190e-03, -6.0375e-03,  5.2883e-03, -1.6542e-03,
         -4.5450e-03, -1.8576e-02, -6.1301e-02,  1.1251e-02, -1.4227e-03,
          1.9841e-02,  3.2629e-02, -3.8623e-02,  4.3724e-02,  2.8845e-03,
         -1.2623e-03, -3.3896e-02, -3.3633e-02,  7.1120e-02, -2.6030e-03,
         -2.8297e-03, -8.0999e-03, -4.7974e-02,  4.8721e-02, -1.7168e-02,
          1.9539e-02, -2.5681e-03, -1.0760e-02, -1.8923e-02, -3.6681e-02,
          4.5460e-02, -3.8324e-03, -2.4408e-03, -4.6963e-03, -6.3194e-02,
          4.6250e-02, -2.0569e-03, -6.8971e-02, -1.2619e-02, -1.3678e-02,
          2.7643e-03, -5.0368e-02,  4.6369e-02, -7.0448e-02, -4.9658e-02,
          2.0162e-03, -1.9849e-02, -3.8212e-02,  2.5966e-02,  5.9269e-03,
         -2.2679e-03,  2.7198e-02, -1.6954e-02,  8.4368e-02, -5.9177e-02,
          3.0999e-02,  3.8469e-02, -7.1604e-02, -5.3525e-02, -2.4468e-02,
         -3.6728e-06,  3.3079e-02, -7.7069e-02, -6.8721e-02,  4.9685e-02},
        '{ 8.2576e-02, -1.3214e-02, -4.2874e-02,  1.4542e-01,  1.0391e-01,
          1.0991e-01, -1.0615e-03, -4.1736e-02,  6.2445e-02,  1.4691e-01,
          2.5425e-02, -1.0696e-01, -1.9330e-02, -6.3385e-02, -3.2138e-02,
         -1.1070e-01,  2.7039e-02,  7.5285e-02, -1.0888e-01, -1.3418e-01,
         -4.8438e-02,  7.0497e-02,  1.6163e-01,  1.2542e-01,  4.0775e-02,
         -3.8326e-02,  5.0664e-02,  7.7969e-02, -1.9080e-02, -1.2172e-01,
         -2.2881e-03, -1.0094e-01, -1.6751e-01, -4.6707e-02,  1.8024e-03,
         -1.8325e-01, -5.9631e-02,  1.3302e-01,  1.4853e-01, -8.5887e-02,
          9.5133e-02, -8.8353e-02,  4.3619e-02,  5.7195e-02, -1.7839e-02,
          5.5511e-02,  2.1413e-02, -1.3435e-01, -1.3275e-01,  1.3711e-01,
         -3.8721e-02, -9.1203e-02,  1.3090e-01,  8.2930e-02, -1.6421e-01,
         -5.4004e-03,  7.9391e-02,  3.3248e-02, -7.4399e-02,  1.1679e-01,
         -4.8404e-03,  1.0077e-01,  1.2733e-01,  1.2200e-01,  1.3547e-02,
          6.2841e-02, -4.1821e-02, -2.2997e-02,  9.1400e-02, -4.9988e-02,
          5.6393e-02, -1.8325e-01, -7.6050e-02, -1.7892e-01, -5.0383e-02,
         -4.2601e-02, -4.3170e-02, -7.6285e-02, -3.5925e-02, -2.8136e-03,
          1.5894e-02,  1.5935e-03,  7.1931e-02, -1.5587e-02,  4.4107e-02,
          1.8088e-02, -4.2779e-02,  1.0333e-02,  9.7548e-02, -1.2295e-02,
          9.9937e-02,  1.0486e-01, -1.0849e-01,  8.5662e-02,  1.2129e-01,
          3.6441e-03, -1.6752e-01, -5.1278e-02, -4.9959e-02,  7.1629e-02,
         -1.5694e-01,  2.6449e-02,  8.7197e-02, -1.0234e-01, -1.0731e-01,
         -1.7995e-01, -3.9433e-02,  8.9750e-02,  6.4226e-02, -1.4028e-02,
          4.8455e-02, -1.0995e-01, -2.3232e-02, -1.4240e-01,  1.5848e-01,
         -9.2622e-02,  4.3590e-02, -1.9229e-01, -7.2645e-02,  5.4355e-02,
          9.9475e-02,  9.8208e-02,  8.8151e-02, -1.5912e-01, -3.7063e-02,
          1.2943e-01,  2.1385e-02,  1.1730e-01, -4.6127e-02, -3.0235e-02,
          3.8753e-02, -7.4115e-02,  2.1794e-02,  1.0951e-01, -4.5406e-02,
          9.1054e-02, -7.0948e-02,  3.6286e-02,  1.4083e-01,  3.6259e-02,
         -4.2758e-02, -1.1574e-02, -1.0938e-01,  8.9624e-02, -1.8706e-02,
          1.2113e-01,  5.8666e-02, -1.3869e-01, -9.7353e-02, -9.4316e-02,
         -1.6000e-01, -1.5090e-01, -1.5692e-01, -1.2744e-01,  5.0359e-03,
         -1.1012e-01,  1.0014e-01, -9.8434e-02,  6.0241e-02,  1.7560e-02,
          2.4315e-02,  6.9601e-02,  9.8229e-02, -8.7925e-02, -8.9978e-03,
          7.2962e-02,  6.2969e-02, -1.7157e-01,  6.7494e-03, -1.0358e-02,
          5.9382e-03,  7.3589e-02,  5.9436e-02, -4.9465e-02, -1.0048e-01,
         -1.6363e-01, -2.3118e-02, -1.2182e-01, -1.1636e-01, -7.1248e-02,
         -1.0514e-01,  2.7379e-02,  1.3876e-01,  1.3425e-01, -2.0220e-02,
          1.0100e-01,  1.4485e-01, -8.2639e-02,  1.1184e-02,  5.0909e-02,
          1.6588e-01,  1.2580e-01, -8.0390e-03, -5.0381e-02,  1.2490e-01,
         -9.5660e-02, -1.3032e-01, -1.0135e-01, -6.9281e-02,  1.2264e-02},
        '{-1.1184e-01,  1.1740e-01,  1.8915e-01,  1.5376e-02,  1.6435e-01,
          1.3910e-01,  9.8743e-02, -5.0672e-02,  1.2707e-01,  8.9991e-02,
         -4.0806e-02,  8.8057e-02,  1.2345e-02, -1.5157e-01, -7.2764e-02,
         -2.3805e-02,  6.9999e-02,  5.7238e-02,  1.3838e-02,  1.2318e-01,
          5.5336e-02, -1.1529e-01, -5.4215e-02, -1.6101e-01, -5.0127e-02,
          5.3783e-02,  2.6618e-01,  1.2019e-02, -1.0145e-01, -9.9731e-02,
          2.8927e-01,  5.6694e-02,  2.8010e-01,  1.3753e-01, -2.1543e-01,
          1.2422e-01,  9.5535e-02,  1.9847e-01,  5.7557e-02,  5.9951e-02,
          3.2160e-02,  1.0314e-01,  1.8910e-02, -1.5667e-01,  2.7720e-01,
         -1.6752e-01, -1.4597e-01, -2.7109e-02, -1.1963e-01,  1.9110e-01,
          2.6219e-02, -3.3848e-02, -1.5491e-01, -3.4467e-02, -6.8710e-02,
         -1.4394e-01,  5.0259e-02,  1.5142e-01,  1.3872e-01, -1.9529e-02,
          2.3601e-03, -1.1315e-01,  1.1591e-01,  1.3299e-01, -5.0143e-02,
          6.9228e-02, -1.6327e-01, -1.3559e-01, -8.1905e-02, -3.7262e-02,
         -8.3456e-02,  2.0561e-02,  2.7204e-02, -8.7203e-02,  6.9294e-02,
         -8.9670e-02, -1.2017e-01, -1.9763e-01, -1.6279e-01, -1.9134e-01,
         -7.9126e-02,  1.6167e-02,  4.8388e-02, -1.3286e-01, -9.8649e-03,
         -1.2241e-01,  1.4059e-02, -2.5653e-02, -3.2184e-02,  1.2793e-01,
         -7.0029e-02, -1.1293e-02,  7.2778e-02,  1.0841e-01, -1.0760e-01,
         -8.0609e-02,  1.4164e-01,  3.1059e-02, -1.1493e-01, -2.4597e-01,
          7.3617e-02,  1.0343e-01,  1.9846e-03,  1.1144e-01, -9.0902e-02,
          1.2876e-01, -1.6903e-02,  1.2783e-01, -3.1852e-03,  7.1692e-02,
          7.5723e-03,  3.8400e-02, -1.0924e-01,  8.1618e-02, -1.4129e-02,
          5.2899e-02,  2.7667e-02, -5.4705e-02, -1.2914e-01, -3.4016e-03,
          2.1842e-03, -1.2408e-01,  1.1452e-01,  5.0309e-02, -1.2590e-01,
          8.6310e-02,  1.2706e-01,  1.8711e-01,  1.4607e-01, -1.0854e-01,
          4.1344e-02,  2.6706e-01,  2.8753e-01,  2.8496e-01,  2.4907e-02,
          5.6483e-02,  6.2425e-02, -1.5850e-01, -1.0077e-02, -8.8933e-02,
         -9.6315e-02, -1.0774e-01,  2.7355e-02,  1.0200e-02, -2.3215e-02,
          2.9433e-02,  3.3507e-02, -1.0142e-02,  2.5949e-02,  1.5768e-01,
         -4.9475e-02,  7.9289e-02, -9.4605e-02, -3.1927e-02,  6.3590e-02,
          1.2259e-01, -5.5264e-02,  1.3314e-01, -6.6328e-02, -2.5635e-02,
         -1.4380e-01,  1.2689e-02, -1.6818e-01, -5.3818e-02,  2.2764e-02,
          8.8323e-02,  4.5771e-02, -1.9549e-02,  1.7838e-01, -7.6911e-02,
          4.7799e-02,  1.0974e-01,  1.2366e-02, -2.5396e-02, -8.4059e-02,
          1.4348e-02,  9.0699e-02, -7.6509e-02,  1.2526e-01,  8.9412e-02,
          1.6357e-02, -2.7005e-02,  1.3307e-01, -8.5769e-02, -2.9203e-02,
          1.2798e-01, -7.6126e-03, -2.1007e-02,  3.6718e-02,  1.0228e-01,
          1.0115e-01,  1.3673e-01, -1.5028e-01,  9.0609e-02, -6.9354e-02,
          5.8244e-02,  5.8260e-02, -1.5317e-01,  3.9882e-02, -1.3967e-01},
        '{ 8.2934e-04, -9.1079e-02,  3.1208e-02,  1.4767e-01, -1.1235e-01,
          6.8007e-02,  5.9675e-02,  9.1962e-02,  1.7301e-01,  4.0595e-02,
          5.1090e-02,  8.3826e-02, -1.7370e-01, -1.9521e-02,  1.0390e-01,
         -6.0303e-02, -4.7017e-02,  1.1589e-01,  3.1827e-02,  9.1108e-02,
         -1.2910e-02, -6.4818e-02, -2.2047e-01,  1.1676e-01, -7.7671e-02,
          1.3949e-01, -7.7835e-03,  3.7735e-02, -1.4179e-01,  7.1374e-02,
          1.3615e-01,  2.4686e-01,  8.8481e-02, -3.0890e-01, -9.7388e-02,
          3.9514e-02,  6.6491e-02,  1.2452e-01,  6.6453e-02, -6.2392e-02,
          1.4222e-02,  9.8804e-02,  1.9197e-01,  7.6411e-02, -5.5808e-02,
          9.1253e-02,  1.8089e-01,  3.1823e-02,  9.0572e-02, -2.5823e-02,
          6.6154e-02, -4.5672e-02,  6.0072e-02,  3.0067e-01,  9.6979e-02,
         -2.4487e-02,  1.0653e-01,  2.1112e-01,  2.0491e-03, -4.5096e-02,
          1.7920e-01, -1.0880e-01,  1.3874e-01,  1.6832e-01, -1.4422e-01,
          1.4820e-01,  2.6271e-02, -7.6557e-02,  4.2831e-02, -1.1337e-01,
          3.3740e-02, -4.5856e-02,  8.1357e-03,  1.0488e-01,  2.1438e-01,
         -2.3265e-02, -4.0760e-02, -2.5522e-02,  9.9530e-02,  1.3467e-01,
          8.3716e-02,  7.3391e-02,  1.2567e-01,  9.1409e-02,  8.1709e-02,
         -4.8238e-03, -1.1831e-01,  9.8311e-02,  2.9682e-01, -7.9560e-02,
         -6.0465e-02,  7.2772e-02,  9.4885e-02,  7.5424e-02,  4.7790e-02,
         -8.6377e-02, -3.7866e-02,  1.4824e-01,  8.2939e-02,  7.1528e-02,
          9.7402e-02, -3.4774e-02, -9.5808e-02, -6.8261e-02, -8.2849e-02,
          1.2402e-01,  3.2234e-02,  9.1089e-02,  2.3137e-02,  4.0195e-02,
         -2.2505e-02, -1.3853e-01, -5.5095e-02, -4.6310e-02, -1.1337e-01,
          6.7064e-02, -8.3180e-02,  1.3578e-01,  1.7633e-02, -1.0262e-01,
         -1.6141e-01, -2.2964e-02,  1.0649e-01,  1.3116e-01, -1.3491e-01,
         -1.4470e-02,  1.1119e-01,  5.7015e-02, -2.3770e-01, -1.6287e-01,
         -3.9919e-02,  3.0985e-03, -1.8277e-02, -3.3250e-02, -1.1710e-01,
         -3.4296e-02, -1.8500e-01, -5.2772e-02,  1.1757e-01, -2.9461e-02,
          1.1043e-01,  1.3280e-02,  5.7240e-03,  1.4476e-01,  5.3430e-02,
          6.6571e-02, -1.0541e-01,  1.4900e-01,  1.8662e-01, -7.5955e-02,
         -1.3947e-01, -1.1089e-01, -1.4791e-01,  1.7765e-01,  5.5108e-02,
          4.4763e-02, -1.6006e-02,  9.3355e-02, -1.2727e-02,  8.7621e-03,
          1.0741e-02, -5.9649e-02,  1.1304e-01,  2.3197e-01, -1.0313e-01,
          1.1738e-01, -1.1260e-01, -4.6185e-02,  1.2053e-01, -1.2115e-01,
          2.4797e-02,  5.0465e-02, -9.7093e-02, -5.8345e-02, -9.3760e-02,
          5.0697e-02, -5.2428e-02,  7.6215e-02,  6.0156e-02, -6.3922e-02,
         -7.3827e-02, -1.0191e-01,  9.4294e-02,  5.1136e-02,  7.9326e-02,
          3.3949e-03, -1.2427e-01,  1.7610e-02,  1.9875e-01,  5.4646e-02,
          1.1426e-01, -1.5676e-01,  6.1511e-02,  3.9180e-03, -1.3031e-01,
         -3.2578e-02,  5.6153e-02,  3.7131e-02,  9.7810e-02,  8.2596e-02},
        '{-6.2647e-02,  6.9348e-02,  4.8825e-02,  8.2631e-02, -1.7519e-02,
          2.2913e-03,  1.5845e-02, -9.5469e-02,  9.0002e-02,  1.3824e-02,
          7.0787e-03, -5.2917e-03, -2.4157e-02,  2.5095e-02, -6.1973e-02,
         -2.3335e-03, -7.6810e-03,  3.5140e-02, -4.0274e-04,  3.7721e-02,
         -1.2036e-03,  6.4069e-03, -7.4290e-02,  8.2113e-02, -2.9723e-02,
          5.6832e-03,  1.4737e-04, -1.9829e-04, -3.9238e-03,  1.0827e-02,
          1.0781e-02,  5.0617e-02,  4.0997e-02,  3.0484e-03,  1.4673e-02,
         -8.6862e-03, -6.0025e-03,  5.4237e-02,  1.0682e-02, -7.6646e-03,
          1.4525e-02,  1.1360e-02, -6.4423e-03, -3.9515e-04,  1.4320e-02,
          5.3167e-03,  6.9265e-03, -4.1790e-04, -2.6774e-02,  3.4407e-02,
          1.3096e-02, -1.2234e-02, -1.4278e-03,  1.5771e-04,  5.7175e-04,
         -3.6705e-03,  2.8178e-02,  8.4498e-03, -2.1077e-02, -1.0294e-03,
         -3.3711e-03, -2.5922e-02,  4.9247e-02, -3.8422e-02, -7.9767e-04,
         -4.6075e-03, -8.3590e-04,  1.7646e-02,  4.8250e-02, -5.5368e-03,
         -4.0491e-04, -3.6019e-02, -2.8340e-03,  1.6864e-02,  4.8279e-04,
         -4.7260e-03, -3.3750e-02, -4.7597e-04, -1.4035e-04,  1.5981e-04,
         -1.0595e-03, -4.0037e-02, -8.3215e-03, -7.8421e-03, -7.6660e-05,
         -1.8772e-03, -2.1871e-03, -6.2557e-03,  3.7423e-02, -8.2944e-09,
          1.0028e-04,  2.8653e-05,  7.6849e-03,  2.0753e-02,  1.9928e-05,
         -8.1122e-05, -1.3439e-02, -8.8735e-03, -3.3653e-02,  4.8218e-06,
          3.8279e-02, -8.7456e-02, -5.0688e-02, -5.0412e-02,  3.0567e-03,
         -4.8067e-02,  7.5471e-02, -7.7559e-02, -6.8093e-02,  3.1730e-02,
         -6.8699e-03, -9.5858e-03,  1.7855e-02,  1.9055e-03, -2.5960e-02,
          9.8089e-04, -5.8628e-04, -6.7784e-02,  3.6670e-03, -6.9661e-02,
         -4.0255e-04,  5.4247e-03,  7.2637e-02, -4.9525e-02, -1.2054e-02,
         -3.2194e-03, -3.4617e-03,  1.2552e-03, -2.5992e-05, -1.9356e-03,
          7.1707e-03,  5.6499e-02,  2.1569e-02, -3.9812e-02, -5.4273e-04,
         -1.7153e-03, -2.0553e-02,  1.1478e-02,  4.3990e-02,  1.9021e-02,
          1.4403e-03, -6.1095e-04, -2.4486e-02,  7.4729e-03, -2.7311e-03,
         -6.1648e-04, -1.0310e-03, -4.0136e-03, -4.0345e-02, -2.6384e-02,
          4.1489e-03,  6.8714e-02, -4.0955e-03, -3.5908e-03, -9.1754e-03,
         -1.1840e-02,  3.6702e-02, -4.2621e-02,  8.9509e-02, -4.2898e-02,
         -4.7971e-03, -2.0877e-03, -5.8819e-02, -4.9264e-03,  5.0281e-02,
         -2.4783e-03, -1.6486e-04, -6.8880e-02,  1.0284e-01, -5.4321e-02,
         -3.1458e-04,  5.9136e-03,  4.6079e-02, -2.2821e-02, -4.3008e-02,
          4.3811e-02, -4.2090e-02, -6.3361e-02, -7.3156e-02, -1.4472e-02,
          6.9004e-03,  2.2154e-02,  8.3692e-02,  5.0320e-02, -1.5502e-02,
         -8.5859e-03, -9.2853e-03, -9.4978e-02, -9.7420e-02, -8.0568e-02,
         -8.6232e-04, -1.1435e-03, -4.1489e-02, -8.3538e-02, -7.2266e-02,
         -1.3482e-03, -5.1673e-03,  1.6240e-03, -5.8643e-02, -7.0320e-02},
        '{ 3.3974e-02, -2.7523e-02,  1.8352e-01, -5.5113e-02,  4.7951e-02,
          1.1836e-01,  6.1956e-03, -4.4113e-02,  1.6972e-01,  2.0955e-02,
          1.0213e-01, -6.5734e-02, -1.3376e-01, -1.7962e-01, -1.1494e-01,
          3.1537e-02,  1.7863e-01,  9.0714e-02, -3.5513e-02, -8.7561e-03,
          7.0112e-02,  1.2929e-01, -2.0643e-01, -9.1320e-02, -1.1601e-01,
          2.4976e-02, -8.1211e-02,  7.9233e-02,  3.4105e-02, -1.4313e-01,
         -6.4392e-02,  1.9517e-01,  8.4059e-02, -7.6107e-02, -1.2814e-01,
         -1.5988e-02,  1.2623e-01,  1.4550e-01, -9.4676e-03,  4.6484e-02,
         -2.5462e-02,  9.1655e-02,  2.1854e-01, -1.0644e-01,  2.8759e-02,
          5.1958e-02,  6.8688e-02,  7.1199e-02, -6.1578e-02, -1.6084e-01,
         -4.2844e-02, -1.4373e-01, -1.8761e-02, -1.2524e-01, -8.3311e-02,
          4.6454e-03,  1.7249e-02,  8.5995e-02,  7.0685e-02, -1.9210e-02,
          7.7310e-02,  6.1377e-02,  2.7909e-04,  2.2946e-01, -4.8738e-02,
         -1.2117e-01,  1.2240e-01,  1.4717e-01,  1.2071e-01, -1.5727e-01,
         -1.4212e-02,  8.9840e-02, -2.1247e-02,  1.2226e-02, -3.5558e-02,
         -1.3004e-01, -4.0356e-02, -9.9225e-03, -2.1706e-02, -1.1384e-01,
          4.8450e-02,  1.6491e-02, -1.0446e-01,  3.2300e-02, -4.4966e-02,
         -1.4421e-01,  7.4976e-02, -8.9343e-02,  1.1276e-02, -7.2893e-03,
         -8.6801e-02,  6.2377e-02, -2.9969e-02,  2.5487e-01,  7.8740e-03,
          5.5174e-02,  4.9402e-02,  1.7232e-01,  1.2369e-01,  5.7131e-03,
         -1.0566e-01, -1.5359e-01,  6.1127e-02, -7.6563e-02,  1.0009e-01,
         -1.1620e-01,  1.4153e-01, -4.9274e-03,  2.2922e-01, -6.0599e-02,
          6.3522e-03,  7.5588e-02, -1.1912e-01,  8.0968e-03,  2.1576e-02,
         -5.4818e-02, -1.5543e-01, -2.0573e-01,  1.2184e-01, -9.4990e-02,
          1.2361e-01, -2.8922e-02, -3.5195e-02,  7.0157e-02,  4.1225e-02,
         -4.5770e-03, -1.2420e-01, -2.5751e-02, -2.0129e-01, -1.5029e-01,
          1.0794e-01,  4.3956e-02,  2.2524e-01,  1.6518e-01,  8.5684e-02,
         -9.1769e-02,  6.7549e-02,  1.3191e-01,  1.0321e-01, -1.1877e-01,
          2.1946e-01,  6.0059e-02,  1.2294e-01,  1.4015e-01,  4.6718e-02,
         -2.4388e-03, -2.0826e-01, -4.0448e-02,  3.5847e-02, -4.7810e-02,
          1.2623e-01,  7.9054e-02,  1.0714e-01, -1.2474e-01,  1.0011e-01,
         -4.1896e-02,  1.4307e-01,  1.4884e-01, -3.6516e-03,  1.4673e-01,
         -8.6925e-02, -6.9808e-03, -4.2107e-02, -1.4266e-01, -8.2891e-02,
         -1.2566e-01,  8.2231e-02, -8.1450e-02, -3.3589e-02,  1.2543e-02,
          1.0368e-01, -8.8106e-02,  9.1006e-02, -1.2165e-02, -1.8446e-01,
         -6.3149e-02,  4.0279e-02, -3.9026e-02,  5.6916e-02,  1.4896e-02,
         -5.7563e-02, -3.9010e-02,  8.6065e-02,  1.3522e-01,  5.1556e-02,
          2.1716e-02,  7.3428e-02, -7.0848e-02,  4.9862e-02,  8.1798e-02,
          1.2849e-01, -3.2286e-02, -1.3132e-01, -7.8957e-02,  1.2871e-01,
         -9.8238e-02,  2.1380e-04,  5.4968e-02, -1.4425e-01, -1.7762e-01},
        '{ 3.5423e-02,  2.8908e-03, -1.3516e-02,  7.3615e-02,  1.3440e-02,
          7.6438e-02, -3.8424e-02, -1.0792e-01,  4.6824e-03, -8.2051e-02,
          3.3059e-02, -3.1193e-02,  1.5704e-01,  2.4905e-01,  2.1048e-01,
         -2.0162e-02, -2.1177e-02,  7.8236e-02, -1.7250e-01,  5.1773e-02,
         -6.9774e-02,  1.3270e-01, -8.1937e-02,  6.2597e-02,  2.1559e-01,
          4.6831e-02,  1.6091e-01,  1.2533e-01,  9.2811e-02,  3.5006e-01,
         -1.7714e-01, -5.9146e-02,  1.5530e-01,  2.3266e-01,  1.4951e-01,
          1.4171e-01, -1.1511e-03,  1.0534e-01,  1.9974e-01,  1.8625e-01,
         -9.8048e-02,  2.1126e-02,  2.2053e-01,  8.8501e-03, -9.7296e-02,
          1.4699e-01,  3.2572e-02,  3.0234e-02,  1.7786e-01, -4.4137e-02,
          1.3016e-01, -8.0046e-02, -1.0226e-01, -1.1250e-01, -1.1813e-01,
          1.4784e-01, -5.9761e-02,  7.3555e-02,  4.2077e-02,  6.5830e-02,
          1.4869e-01,  6.5118e-02, -3.4468e-02, -4.8266e-02, -5.9225e-02,
         -8.0890e-02, -9.3814e-02, -1.1015e-02, -3.2928e-02, -4.3897e-02,
          4.8567e-02,  4.8863e-02, -1.6283e-01,  1.1889e-01,  2.2105e-02,
         -5.2072e-02, -1.0028e-01, -4.8980e-02, -1.6344e-01, -2.3617e-01,
          4.3386e-02,  9.5878e-02, -1.3813e-01, -1.1958e-01, -1.4034e-01,
          1.3681e-01, -9.0166e-02,  4.8030e-02, -9.2500e-02, -1.0783e-01,
         -7.1062e-02, -1.6627e-01, -1.6373e-01, -1.4834e-01, -2.2686e-02,
          6.7022e-02, -5.9591e-02, -6.9549e-02, -2.9621e-02, -1.4252e-02,
         -4.8838e-02,  7.6882e-02,  1.9600e-01, -6.3742e-02,  3.8135e-02,
         -7.9644e-04, -4.4097e-02,  6.9348e-02, -1.0155e-01,  8.4934e-02,
         -1.2192e-01,  8.1246e-03,  1.3737e-02,  6.4013e-02, -7.8701e-02,
          6.7624e-02,  4.7999e-02,  1.6201e-01,  7.7419e-02,  1.3040e-01,
         -8.8261e-02,  6.3101e-02,  1.2149e-01,  1.0504e-01,  6.3741e-02,
          3.1296e-02,  3.0441e-02,  1.2541e-01,  9.8311e-02,  2.0964e-01,
         -7.5340e-02,  1.8893e-01,  1.2297e-01,  1.4246e-01,  1.3420e-01,
          2.9589e-02,  3.1539e-03, -7.3998e-03, -7.5072e-02,  8.6288e-02,
          2.9794e-02,  1.6061e-01,  3.0367e-02,  1.2790e-01, -7.4691e-02,
          1.0141e-01, -4.2026e-02,  1.2555e-01, -5.4209e-02,  4.3931e-02,
          6.8367e-03,  8.3907e-02, -7.7789e-02,  1.6579e-01,  7.5851e-02,
         -8.5639e-02,  9.7931e-02,  1.3363e-01,  7.7576e-02,  2.5825e-02,
          4.1565e-02,  7.3223e-02, -1.1416e-01,  9.2078e-03, -5.6158e-02,
          7.5485e-02,  8.2947e-02,  1.6436e-01, -5.7661e-02, -1.1858e-01,
          1.7586e-01, -3.8256e-02,  1.0953e-01,  5.3639e-02, -4.1900e-02,
          2.9562e-02, -5.4470e-02,  1.2995e-01, -5.0640e-02, -9.7492e-02,
         -4.8673e-02,  2.0655e-02, -6.7979e-02, -1.4128e-01, -8.0460e-02,
         -1.2362e-01, -3.4179e-02,  7.3192e-02,  2.2818e-02, -2.5338e-02,
          1.8109e-02,  4.2519e-03,  1.4896e-01, -7.7530e-02, -9.5053e-02,
          1.4282e-01, -8.0049e-02,  7.7640e-02, -8.7395e-02,  1.9694e-01},
        '{-6.8487e-02, -5.0296e-02,  1.3742e-01, -1.5139e-01, -1.2365e-01,
          1.7622e-02, -4.8330e-03, -1.1720e-01, -1.7492e-04,  1.0532e-01,
         -6.1933e-02,  3.4548e-02,  5.0355e-02, -3.7451e-02,  7.7647e-02,
         -5.3012e-02,  2.8783e-02,  7.9195e-03,  1.6259e-01, -6.1120e-02,
          1.7994e-01,  1.3471e-01,  2.5976e-01, -6.8551e-02,  3.7579e-02,
         -1.2384e-01, -5.1189e-02,  9.6477e-02, -5.6043e-02,  1.1652e-01,
         -4.0215e-02,  1.2083e-01,  3.6784e-02,  5.0062e-02,  1.9949e-02,
         -2.8896e-02, -1.3837e-01, -8.6966e-02,  2.3010e-01, -1.0338e-01,
         -2.7594e-02,  1.0905e-01,  1.5743e-01,  9.8341e-02, -1.8406e-01,
          7.1670e-02,  4.7352e-03,  5.2448e-02,  2.0577e-01,  9.5951e-02,
         -2.6488e-02, -1.1093e-01, -1.2710e-01, -1.5263e-01,  2.9924e-02,
         -1.0604e-01,  2.0949e-02,  5.1720e-02, -5.8880e-02,  3.2519e-03,
         -1.2285e-01,  9.2454e-02, -3.1067e-02,  8.0896e-02,  5.9996e-02,
         -7.3132e-02,  4.1940e-03, -1.4423e-02,  3.6550e-02, -9.6402e-03,
         -1.4427e-01, -9.5249e-02,  4.2483e-02, -1.5881e-01,  4.4422e-02,
          7.7040e-02, -8.4667e-02, -6.5250e-02,  5.8374e-02,  1.4803e-02,
          6.1323e-02, -8.9839e-02, -1.0727e-01, -2.9680e-02, -1.3307e-01,
          2.2125e-02, -4.9086e-02,  1.5598e-01,  3.5020e-02, -1.0565e-01,
          1.7012e-02,  1.1895e-01, -1.8501e-01, -1.2878e-01,  1.2353e-01,
         -5.4019e-02,  5.3103e-02, -5.6720e-02, -3.6364e-03, -6.7203e-03,
          1.6123e-01,  1.4045e-01,  1.6894e-03,  3.9255e-02,  9.3369e-02,
         -1.0621e-02, -1.7489e-01,  8.7540e-03,  1.5720e-01, -1.7668e-01,
         -1.7309e-01,  7.0994e-02,  4.0360e-02, -2.0236e-01,  9.5876e-02,
         -1.3067e-01, -2.6941e-02, -1.8481e-01,  5.6618e-02,  1.7502e-01,
          1.5670e-01,  4.2189e-02,  1.1566e-01,  7.9337e-02,  1.7811e-01,
          3.8871e-02,  6.6160e-02,  1.8489e-01, -1.1374e-01, -1.0067e-01,
          5.5282e-02, -7.3313e-02, -3.2874e-02, -4.6636e-02,  1.5365e-01,
          2.8468e-02, -9.1009e-02, -4.0409e-02,  1.7941e-02,  3.4543e-02,
         -1.6288e-01,  1.4257e-01,  1.4741e-02, -1.7999e-01, -4.8616e-02,
          2.6831e-02, -5.1253e-03, -3.5793e-02, -1.9124e-02,  8.2461e-02,
         -3.1115e-02,  1.1747e-01,  3.9199e-02,  9.6136e-02, -1.5183e-01,
         -4.9133e-02,  5.8133e-02, -8.8241e-02,  1.5122e-01, -1.1437e-01,
          1.0690e-01,  1.5407e-01, -3.0953e-02,  2.8057e-02,  3.6063e-02,
         -7.2424e-02,  4.8382e-02,  4.4845e-02, -1.0202e-02,  9.5907e-02,
          1.3264e-02,  3.3215e-02,  1.7227e-01,  4.5636e-02, -5.8589e-02,
          2.1612e-02,  1.3323e-01, -1.0725e-02, -1.0558e-01,  1.0457e-01,
         -2.9483e-02, -1.6460e-01,  2.7685e-02,  1.4044e-01, -9.4184e-02,
          4.9204e-03,  1.9177e-03,  2.5936e-02, -9.7414e-02,  5.5610e-02,
          6.6316e-02,  3.0586e-02, -1.1390e-01, -4.8380e-02,  6.5991e-02,
         -2.7872e-02, -6.0194e-02, -5.8273e-02, -2.3191e-02,  2.7089e-02},
        '{ 1.2194e-01,  1.1605e-01, -6.2620e-02, -8.1474e-03, -1.5487e-01,
          6.8588e-02,  1.3455e-01,  3.8509e-02,  9.3612e-02,  1.2170e-01,
         -3.3852e-02,  1.2305e-01, -1.4034e-01,  5.4082e-02,  1.1663e-01,
          2.1039e-02, -3.2202e-02,  3.3412e-02,  2.4727e-02,  6.7533e-02,
          1.8078e-01,  8.6966e-02, -4.1365e-02, -1.6803e-01,  9.8777e-03,
         -8.5941e-02,  1.4568e-01,  1.0989e-01,  4.2275e-02, -4.1596e-02,
          7.5711e-02,  4.9881e-02,  6.2601e-02, -4.0431e-02, -1.2012e-01,
         -2.8566e-02,  3.0408e-02,  2.3573e-03, -6.8083e-02, -1.5128e-01,
          1.2339e-01, -1.0811e-02,  7.7769e-02, -9.6633e-02, -4.6987e-02,
         -1.2676e-01,  3.6679e-02,  6.7116e-02,  3.8837e-02,  1.7290e-01,
         -2.4725e-02, -7.0026e-02, -2.2962e-02,  7.5442e-02,  8.0203e-02,
          9.2967e-02, -2.0109e-02, -1.0908e-02, -1.3480e-02, -4.5244e-02,
         -7.1990e-02, -1.8520e-02,  1.1060e-01,  6.5080e-02, -1.4334e-01,
          1.1260e-02,  5.9300e-02, -1.4951e-01, -2.3908e-02,  2.8395e-02,
         -3.4244e-02,  4.9056e-02,  6.6137e-02, -1.1482e-02, -1.3091e-01,
         -1.0511e-01,  8.8006e-02,  7.8426e-02,  6.0506e-02, -6.3731e-02,
          1.1525e-02,  2.2355e-02,  8.3377e-02,  2.8695e-02, -4.4691e-02,
         -1.1082e-01,  3.5650e-02,  8.3314e-03,  5.9749e-02,  1.0820e-01,
          6.4583e-02,  7.7160e-04,  7.7803e-02, -9.2524e-03,  1.8444e-01,
          2.7806e-02, -4.5384e-02,  9.1867e-02,  4.2767e-03, -7.1033e-02,
         -1.2864e-02, -3.3713e-02, -7.3554e-02,  1.1643e-01, -1.8411e-03,
          6.7903e-03, -1.1577e-02, -1.0943e-01,  9.8626e-02,  2.1052e-02,
          9.7484e-02,  3.9055e-02, -1.1624e-03, -1.1654e-01, -6.2956e-03,
          8.3171e-02, -1.5413e-01,  1.0457e-01, -1.4626e-01, -1.9342e-03,
          1.0483e-02,  2.5168e-02,  6.6272e-02, -1.3429e-01, -1.0167e-01,
          1.1523e-01,  9.1384e-02,  7.9335e-03, -1.6923e-01,  1.8517e-02,
          2.8150e-02,  1.3665e-01,  9.5702e-02, -9.7238e-02, -1.5557e-01,
          3.6423e-02, -9.6864e-02,  7.2188e-02,  9.6425e-02, -8.7708e-02,
          1.5004e-01, -5.4294e-02, -6.6647e-02, -8.4892e-02,  2.2071e-02,
         -1.0036e-01,  7.5585e-02,  1.0067e-01,  6.7508e-03, -5.8903e-02,
         -7.0386e-02,  2.0453e-02, -1.2770e-01,  1.5488e-01, -8.9259e-02,
         -2.5916e-02, -7.5594e-02, -7.8557e-02,  1.8972e-01,  1.1429e-01,
          1.9329e-02, -1.3637e-01,  9.9563e-02,  4.9154e-02,  5.4947e-04,
          5.7791e-02, -7.7256e-02, -4.4807e-02,  7.7387e-02,  1.8314e-01,
          3.3819e-02, -1.3327e-03,  7.4620e-02,  4.6291e-02, -1.3885e-01,
          8.6140e-02, -8.3485e-02, -3.5988e-02,  8.8968e-02, -2.5188e-02,
          2.7915e-02,  5.6842e-02,  1.1966e-01,  1.1239e-01,  1.3550e-02,
         -9.8130e-02, -2.4170e-02,  1.1213e-02,  2.2276e-02, -6.4039e-02,
         -1.1767e-01, -1.0938e-01, -6.5569e-02, -1.3172e-02, -8.0638e-02,
          9.2300e-02, -1.4571e-01,  8.2418e-02, -1.0637e-03, -1.2166e-01},
        '{ 1.6911e-01, -1.4626e-01,  6.5732e-02, -1.7506e-01,  1.3837e-02,
         -7.9398e-02, -8.3971e-02, -6.5905e-02,  1.4714e-01,  7.6090e-02,
          2.8854e-02,  1.6283e-01, -2.0172e-01, -1.7296e-01,  1.1092e-01,
          3.4354e-02,  1.2273e-01,  9.6714e-02,  1.5357e-01,  1.9924e-01,
          2.3646e-01,  5.3149e-02,  1.0058e-01, -1.0631e-01,  1.4685e-02,
         -9.8871e-02,  1.2998e-01,  1.5458e-01,  1.7994e-01,  2.4519e-02,
          1.7694e-01,  2.2938e-01,  1.4227e-01, -1.7615e-01,  1.0546e-02,
          6.2670e-02,  4.0040e-02,  4.3946e-02,  1.5422e-01, -2.3387e-01,
          1.2056e-01,  2.0797e-01, -2.1515e-02, -2.7007e-02,  2.9457e-02,
          1.2480e-01, -2.9470e-02,  2.8814e-01,  9.1505e-02, -3.3137e-02,
          2.4812e-02, -2.9919e-05,  5.5918e-02,  1.9770e-01,  1.7101e-01,
          2.4929e-02,  7.3764e-02, -2.6293e-02, -1.2788e-01, -1.3939e-01,
         -5.3964e-02, -1.0015e-03,  3.5140e-03,  9.8109e-02, -1.3210e-01,
          6.8001e-02, -1.1852e-01,  7.3168e-02, -1.4859e-01,  9.0289e-02,
          4.2427e-02, -7.6337e-03,  5.0605e-02, -4.3622e-02,  1.5779e-02,
         -8.7326e-02,  1.0184e-01,  8.0786e-02,  1.4641e-01,  1.7502e-01,
          5.3175e-02, -1.0583e-01, -1.0807e-02,  2.8318e-01,  5.1523e-02,
         -1.2858e-01,  1.2582e-02,  1.0739e-02,  2.1621e-01, -1.6348e-01,
         -2.6427e-02,  7.9860e-02,  1.0838e-01, -4.3937e-02, -1.3597e-01,
          7.0948e-02, -4.7180e-02,  1.2999e-01, -1.6572e-01, -1.9028e-01,
         -3.9647e-02,  8.2683e-03,  6.1405e-02, -2.7122e-02,  6.4165e-02,
          4.7630e-02,  4.6474e-03, -7.8652e-02,  2.0695e-02, -1.2723e-01,
         -1.5746e-01, -1.6284e-01,  3.7076e-02, -5.6387e-02,  6.1013e-03,
         -1.1144e-01, -9.1367e-03, -8.0329e-02,  1.1347e-01,  7.1394e-02,
         -7.6480e-02, -1.3224e-01,  1.1916e-02,  4.4499e-02,  4.0416e-02,
          1.8347e-01,  2.4924e-01, -4.3530e-02, -6.3367e-02, -7.4647e-02,
          3.1901e-02,  8.3478e-02, -4.1961e-02,  8.7232e-03,  6.0550e-03,
         -6.5490e-02, -1.7685e-01, -1.4281e-01,  1.9644e-02, -1.0686e-01,
          2.2515e-02, -8.5833e-02, -7.5894e-02, -1.2005e-01,  1.8762e-01,
         -1.0720e-01,  2.8914e-02,  9.6117e-02,  1.0372e-01, -7.8185e-02,
          1.3605e-01, -1.2931e-01, -6.8996e-02,  1.0581e-01, -1.1036e-01,
          4.6765e-02, -4.3251e-02,  3.9042e-02,  4.2334e-02, -1.0854e-01,
          2.5297e-02, -1.2076e-01,  9.2376e-02, -6.7018e-02, -1.7001e-01,
         -9.7124e-02, -4.4309e-02, -1.1749e-01, -5.6254e-02,  1.0059e-01,
          1.2808e-01,  6.7739e-02,  1.7261e-01, -1.0098e-01, -1.1003e-01,
          4.7218e-02,  7.0680e-02, -1.5115e-01,  1.1773e-01,  5.8281e-02,
          9.5880e-04, -8.9555e-02, -9.4265e-02,  1.6599e-01, -1.1721e-01,
         -2.8053e-02, -6.5650e-02,  1.3453e-01,  1.3202e-01,  1.2568e-01,
          6.9625e-02,  8.1710e-02,  1.5492e-01,  7.7727e-02,  1.7606e-01,
          7.4972e-02, -1.3089e-01, -7.6740e-02,  3.1373e-02, -1.0359e-01},
        '{ 7.4226e-02,  9.9982e-02,  2.3964e-03, -1.2497e-01,  2.8198e-02,
          4.5592e-02, -1.1464e-01,  1.3305e-02,  5.9745e-03, -1.1273e-02,
          5.1067e-02, -9.0266e-02, -9.4097e-02,  5.8140e-02, -1.0865e-01,
          1.1906e-01,  5.9056e-02, -3.4673e-02, -2.6929e-02,  6.5225e-02,
          1.3280e-01, -1.3679e-01, -6.4118e-02, -8.9340e-03, -1.3028e-01,
         -3.7000e-02, -1.4300e-01, -3.0026e-02, -5.4532e-02,  6.4243e-03,
          1.0328e-01,  7.8270e-02,  1.9263e-01, -8.5719e-02, -3.0415e-02,
          1.5024e-01,  2.4963e-01,  2.0275e-02, -8.2871e-02,  1.7647e-03,
          7.7041e-02,  1.5832e-01,  1.0688e-02,  1.6916e-01,  2.0326e-01,
         -1.0233e-01, -1.3741e-01, -1.5013e-01, -1.7073e-01,  1.5592e-01,
          5.0221e-02, -9.9454e-03,  5.4623e-02,  5.5070e-02,  9.3283e-02,
         -7.5065e-02, -6.5348e-02,  4.7400e-02,  1.3644e-01, -9.5074e-02,
         -1.2304e-01,  1.1871e-01,  1.8731e-01,  1.4739e-01,  2.8038e-02,
          1.3938e-01, -3.0130e-02, -9.4310e-02, -1.5623e-01, -5.4256e-02,
          6.4856e-02,  5.7347e-02,  1.4644e-01,  1.5108e-01,  4.8615e-03,
          7.5347e-02, -7.9810e-02,  2.4769e-02,  9.1026e-02,  1.7782e-01,
          2.8045e-02,  4.7269e-02,  6.6899e-02,  3.4637e-02,  1.7903e-01,
         -1.1474e-01, -5.3276e-02, -2.5537e-02,  9.0004e-04, -1.8364e-02,
         -3.3418e-02, -6.1830e-02,  2.4464e-02,  6.6425e-02, -1.7038e-01,
          1.1025e-01, -7.0729e-04,  5.4887e-02,  4.7867e-02,  2.1845e-02,
         -4.5729e-02, -5.3182e-02, -5.7105e-02,  7.8901e-03, -6.1396e-02,
         -1.1343e-01, -1.2912e-01,  6.6488e-02, -8.3068e-02, -1.0201e-02,
          8.3586e-02, -6.1242e-02,  7.0400e-02, -5.4015e-02,  9.7373e-02,
          1.9281e-02,  6.7171e-02,  1.0386e-01,  7.3737e-02,  7.8349e-02,
          5.2439e-02,  1.0913e-02,  1.3475e-01,  1.4204e-03, -1.4801e-02,
         -1.3211e-02,  2.3266e-01,  1.8407e-01,  8.2313e-02, -6.3069e-02,
          2.0655e-01,  7.3258e-02, -3.1026e-02, -5.7232e-03, -7.6275e-02,
         -4.2573e-02,  6.9853e-02,  1.6736e-02,  7.3756e-02, -1.2847e-01,
          7.4225e-02, -1.4189e-01, -1.0876e-01,  5.9090e-02,  2.1021e-01,
          1.0026e-01,  9.7633e-02, -6.1800e-02, -1.1932e-01, -1.0780e-01,
          8.5167e-02, -6.3378e-02, -5.2864e-02, -1.0064e-01, -9.9485e-02,
          3.4932e-02, -1.6102e-01,  6.9236e-02,  1.2952e-01,  6.5472e-02,
         -4.4082e-02,  7.7104e-02,  1.1023e-01,  7.6546e-02, -3.1600e-02,
          8.3190e-02, -5.3925e-02,  1.4825e-01, -1.2992e-01,  3.3167e-02,
          1.0773e-01,  1.2363e-01,  8.0030e-02, -4.2297e-02, -1.9609e-01,
         -9.3415e-02,  1.6030e-01,  3.6575e-02, -3.1894e-02,  3.7630e-02,
         -1.5759e-01, -1.6767e-01,  8.5946e-02, -2.0527e-03, -1.1887e-01,
          1.4409e-02,  4.6218e-02,  6.8085e-02,  3.5444e-02, -1.0869e-01,
         -3.3294e-02, -1.4057e-01,  9.6744e-02,  1.3367e-01, -1.5097e-01,
          1.7700e-01, -6.9554e-02,  5.4199e-02, -9.9972e-02, -1.9443e-01},
        '{ 4.3111e-02,  9.0785e-03,  1.7894e-01, -8.7130e-02,  1.1815e-02,
         -3.8335e-02,  1.1374e-01,  5.0911e-02,  8.9619e-02,  4.7414e-03,
          5.2295e-02, -1.1817e-02,  1.8194e-02,  8.0887e-02, -4.5481e-02,
          2.3759e-01,  7.1868e-02, -4.4937e-02,  2.6166e-02,  1.5306e-01,
          2.9926e-02,  9.4180e-03,  1.4089e-01,  1.6099e-01,  1.2564e-01,
          1.1901e-01,  5.3369e-02,  9.3687e-03,  5.3982e-02, -1.8552e-01,
          2.4301e-01,  1.7797e-01,  3.3445e-01,  2.5459e-02, -1.9861e-01,
          2.6280e-01,  2.7959e-01,  1.1749e-01,  1.7910e-02,  2.8116e-01,
          1.3467e-01, -2.6665e-02,  1.0753e-01,  5.8074e-03,  7.4161e-03,
         -3.0640e-02, -7.3579e-02, -3.6922e-02,  7.4537e-02,  1.7315e-02,
          9.4755e-02,  4.3681e-02, -1.3841e-01, -4.3195e-02,  1.1800e-01,
          1.4030e-02, -3.9696e-02,  1.2248e-01,  1.0497e-01,  2.1173e-03,
          7.0231e-02,  6.3736e-02, -7.2866e-03,  9.4063e-02, -9.5132e-02,
         -1.6949e-02, -1.7572e-02, -8.2266e-02, -1.7604e-01,  5.5984e-02,
         -3.6513e-02, -2.3419e-01,  4.0037e-02,  1.8242e-03,  2.5950e-02,
         -9.6393e-03, -1.9047e-02, -1.7175e-01, -1.6486e-01, -1.5759e-02,
         -3.3876e-02,  3.7343e-02, -1.5137e-01, -8.9345e-02,  7.7645e-02,
         -2.8084e-02, -1.2226e-01,  5.0450e-02, -3.9654e-02, -1.6451e-01,
          5.4736e-02,  8.0087e-02,  2.6186e-02,  6.3409e-03,  1.8606e-02,
          6.2597e-02, -1.4658e-01,  4.3864e-02, -1.1207e-01,  3.3666e-02,
         -7.4082e-02,  5.1000e-02,  5.4043e-02,  4.9787e-02,  1.0433e-01,
          1.2894e-01, -8.4417e-02,  5.0063e-03,  1.4354e-01,  1.7652e-01,
         -1.1999e-01, -1.2229e-01,  7.6522e-02, -4.9456e-02,  6.4432e-02,
         -3.1005e-02, -6.3023e-02, -1.3207e-01,  1.0389e-01,  6.1580e-02,
          8.1349e-02, -4.0393e-02, -1.1947e-01,  3.3749e-02,  1.6266e-01,
          4.0822e-02,  6.6790e-02,  1.8899e-02,  2.0009e-02, -2.5515e-02,
          1.0855e-01,  3.7484e-02,  3.0403e-01, -9.2579e-03,  1.5222e-01,
         -6.8267e-02,  5.6837e-02,  7.9938e-02,  1.1507e-02,  1.4883e-03,
          9.0885e-02, -3.5736e-02,  1.0931e-01, -6.3357e-02, -3.7613e-02,
          1.1892e-01, -3.9621e-02,  1.4748e-02, -3.9243e-02,  1.0092e-01,
         -9.5769e-02, -3.8690e-03, -8.9136e-04,  1.3371e-01, -1.6097e-02,
          9.2454e-02, -1.4397e-01,  1.1959e-01,  1.7145e-01, -1.1043e-02,
         -9.9024e-02, -6.5889e-02, -2.0818e-02, -4.2416e-02,  5.7016e-03,
          5.2259e-02,  6.2070e-02, -1.4025e-02, -1.4598e-01,  9.2935e-02,
          1.7048e-01,  9.4552e-02,  1.3218e-01, -2.1856e-02,  1.2962e-01,
         -5.6455e-02,  1.1772e-01, -5.2846e-02,  1.6907e-01, -8.4986e-02,
          1.2640e-01, -4.5140e-02, -5.2895e-02,  9.9871e-02, -5.4058e-02,
          1.7299e-02, -1.4325e-01, -5.1168e-02, -1.3840e-02, -7.9861e-02,
          1.0248e-01, -5.7250e-02,  1.2882e-01,  7.4231e-03, -4.3315e-02,
          1.0573e-01, -3.1458e-02, -1.1453e-01, -7.7525e-02, -3.2600e-02},
        '{ 7.1720e-02,  6.7531e-02, -8.8430e-02,  6.8802e-02, -1.3500e-01,
          1.8049e-01, -1.3556e-01, -1.1639e-01,  1.7988e-02,  5.2399e-02,
         -1.2153e-01,  8.7878e-02,  7.2055e-02,  1.0798e-01, -5.1843e-02,
         -7.4274e-02,  6.2624e-03,  1.0531e-02, -7.3590e-02, -2.5303e-02,
         -1.8341e-01, -1.0052e-01,  5.5971e-04,  1.8432e-01, -6.1757e-02,
         -5.0759e-02,  4.8592e-02,  8.2293e-02, -1.3135e-01, -1.0258e-01,
          1.1807e-01, -4.5472e-03, -6.1773e-02, -5.0369e-02,  3.6552e-03,
          1.3441e-01, -1.0713e-01, -6.8303e-02, -1.6498e-01, -1.6057e-01,
         -1.1794e-01, -1.1696e-01,  6.8550e-02, -1.6038e-01,  4.0971e-02,
         -1.8137e-01, -8.0293e-02, -4.7663e-02,  5.9798e-02,  1.6011e-01,
          7.0238e-03, -6.6723e-02,  9.3478e-02, -1.6677e-03,  1.2431e-01,
         -1.3057e-01, -7.0549e-02,  1.6503e-01, -1.1517e-01, -4.9193e-02,
          2.2134e-02, -4.8995e-02,  2.1389e-02, -2.4226e-01, -1.5125e-01,
         -9.1077e-02,  8.6055e-02, -3.2873e-02,  8.8235e-02,  4.9210e-02,
         -1.7747e-01, -8.6723e-02, -6.4784e-02,  1.0854e-01, -7.9778e-02,
         -7.0909e-02,  9.7976e-02, -5.3444e-02,  3.9114e-02,  2.5408e-02,
          3.7427e-02,  7.5224e-02, -4.0705e-02,  2.2638e-02, -2.2694e-03,
          6.3108e-02, -1.1190e-01, -6.8578e-02,  4.7564e-02,  1.3936e-01,
          1.2460e-01,  1.0504e-01,  1.2424e-01, -1.9919e-01,  8.8271e-02,
         -8.2199e-02, -2.9744e-02, -2.1046e-02, -1.1898e-01, -3.9140e-02,
         -1.1041e-01, -5.9690e-02, -2.0703e-02,  2.1721e-01, -6.1255e-02,
         -8.4788e-02, -1.4507e-02,  1.2965e-01,  3.8589e-02, -1.6930e-01,
         -1.3776e-01, -4.5173e-02, -7.9126e-02,  1.3220e-01,  1.2753e-01,
          3.4464e-02,  4.1198e-02, -7.2390e-02,  1.6905e-01,  7.4407e-03,
          6.5930e-03, -9.2589e-02,  9.2601e-02,  1.0704e-01,  1.3330e-01,
          7.8410e-02,  1.3735e-01, -8.4029e-02, -8.9444e-03, -5.5535e-02,
         -1.2455e-01,  4.0036e-02, -1.3658e-01, -7.2269e-02, -1.7082e-02,
          1.3597e-01, -5.6274e-02, -5.7017e-02,  9.8883e-02,  8.6444e-02,
         -5.5104e-02, -7.5163e-02,  6.4864e-02, -8.1118e-02, -1.3405e-01,
          5.8034e-02, -1.1135e-01,  9.0484e-02, -6.1050e-02,  9.9430e-02,
         -1.8599e-03, -1.2383e-01, -1.0802e-02, -1.4116e-02, -1.2398e-01,
          1.2035e-01, -3.5935e-02, -6.4920e-02, -1.0163e-01, -1.4602e-01,
         -6.7011e-02, -1.4567e-01,  1.8491e-01,  2.0770e-01,  2.8974e-02,
          8.7312e-02,  1.0278e-01,  1.0768e-01, -7.5884e-02, -5.9262e-02,
         -3.6861e-02,  8.6706e-02, -3.0814e-03,  7.5927e-02,  1.4318e-02,
          8.5158e-02, -7.6847e-02,  1.2597e-01, -7.6262e-02,  8.1546e-02,
          9.7976e-03,  8.1927e-03,  1.3764e-01,  1.2889e-01, -1.2166e-01,
          1.4724e-03,  8.2344e-03,  7.6536e-02,  2.0153e-01,  4.2094e-02,
          4.3727e-02,  1.4964e-01,  2.1105e-01,  3.1130e-02,  1.2536e-01,
         -1.5072e-01, -9.4469e-02, -6.4312e-02,  1.1520e-01,  1.6179e-01},
        '{-7.9707e-03,  5.0958e-03, -2.5579e-03, -3.1547e-03, -8.9182e-03,
          9.7588e-03, -8.7289e-05, -6.1406e-03, -9.1722e-03, -1.6317e-02,
         -5.1590e-03, -9.6596e-03, -1.0375e-03, -2.7403e-02, -2.2591e-02,
         -1.5671e-02,  6.5890e-04,  2.0494e-03,  7.4020e-02,  2.5137e-03,
         -5.1250e-03, -3.0969e-03, -4.4745e-02, -2.8074e-02,  4.1301e-02,
         -2.4409e-03,  1.4042e-03, -7.9032e-03, -6.0616e-03,  3.0490e-03,
         -5.1304e-03,  3.9510e-03, -1.4036e-02, -7.3142e-04, -9.5900e-03,
         -1.9617e-04, -1.9700e-02, -5.8376e-03, -2.7345e-03, -8.7758e-04,
         -1.7466e-02, -2.7285e-02, -1.2059e-03,  1.1020e-03, -3.3006e-03,
         -4.7146e-03, -3.5810e-03,  7.2225e-03,  2.2147e-03, -5.3185e-03,
          3.6156e-03, -1.7094e-03, -3.5170e-02,  2.2254e-03,  4.0771e-03,
          6.3865e-05, -1.0657e-03, -3.3190e-02,  1.5168e-03, -1.2248e-02,
         -1.4500e-03, -5.9774e-04, -1.3439e-04, -9.4807e-04, -1.3156e-02,
         -1.2270e-03, -6.7106e-03,  2.2351e-02,  1.2896e-03, -1.0741e-02,
         -9.9781e-03, -1.5296e-02, -4.6410e-02,  4.2423e-03, -4.1624e-03,
          4.8511e-03, -1.0879e-03, -3.0887e-03,  1.1334e-03,  2.7001e-03,
          3.1111e-02,  4.8185e-03, -2.7272e-02,  3.1563e-04, -4.3911e-03,
         -1.7279e-03,  1.0591e-03, -3.0727e-02, -4.1287e-03, -7.1149e-03,
         -3.0555e-03,  7.6003e-04,  3.0499e-03, -6.7317e-03, -5.1276e-03,
         -8.8827e-03, -1.4928e-02,  2.0314e-02, -5.8116e-03,  6.8196e-03,
          1.0117e-03, -4.4701e-02, -3.4419e-02, -7.1406e-02, -1.7545e-03,
         -1.3539e-03, -4.1704e-03, -8.3757e-02, -1.0612e-02, -4.3037e-03,
         -2.8716e-03, -5.1802e-03,  2.1390e-02,  1.7135e-02, -5.6294e-03,
         -5.1082e-03, -1.7146e-03,  6.0128e-02, -3.5165e-03, -2.1379e-02,
         -4.2848e-03, -3.2150e-02,  2.5209e-02, -2.7127e-02, -3.6796e-02,
         -3.7227e-03, -4.9729e-03, -2.0825e-03, -5.1581e-03,  3.3682e-03,
         -8.7830e-03, -3.1916e-04, -2.0541e-02,  4.8990e-02, -1.9059e-03,
         -3.3223e-03,  6.6202e-02, -2.3715e-02, -1.0109e-02, -1.6248e-03,
         -5.8943e-03,  6.1469e-04, -5.5537e-02, -6.1783e-03, -4.7028e-03,
         -9.7101e-03, -1.8833e-02,  3.8043e-02, -7.4227e-03, -1.8771e-02,
         -2.9122e-03,  3.4090e-02,  6.0914e-02,  1.0821e-02, -4.5082e-03,
         -5.7353e-02,  6.6703e-02, -5.5277e-02, -2.5867e-03, -2.4559e-02,
          5.1441e-02, -2.4768e-02,  4.0244e-02,  5.3850e-02, -4.6456e-03,
          1.0455e-02, -6.7235e-04, -4.8802e-02, -1.6643e-02,  6.4343e-03,
         -9.3166e-03, -4.8847e-03,  7.7992e-02, -3.8211e-03,  5.0646e-03,
          2.5992e-03,  3.4350e-02,  1.3792e-02,  5.1641e-02,  1.1949e-02,
          3.2063e-02, -4.4037e-03, -3.6912e-03, -4.2405e-03,  4.2587e-03,
          1.0746e-02, -5.1435e-03,  1.5517e-02, -2.7836e-03, -3.3271e-02,
         -8.9573e-03, -1.0165e-03, -6.4922e-02, -4.1450e-03, -1.7512e-03,
         -9.2138e-03, -3.3412e-02, -3.7805e-02, -2.0437e-02, -1.4496e-02},
        '{-7.6217e-02, -9.9469e-02,  9.6388e-02, -1.1528e-01, -1.1294e-02,
          5.0888e-02, -3.2652e-02, -1.8167e-01,  2.7120e-02, -2.5874e-02,
          9.9474e-02, -1.5122e-01,  7.1681e-02, -4.4850e-02,  1.3853e-01,
         -4.2217e-02,  7.7391e-02, -7.6994e-02,  3.5506e-02, -1.1699e-01,
          7.9705e-02, -1.6556e-02,  5.3457e-03,  1.2003e-01, -1.2590e-01,
         -1.2267e-01, -5.8743e-02, -7.6585e-02, -1.0110e-01,  2.4626e-02,
          2.9707e-02,  7.7755e-04, -1.5710e-01, -5.9428e-02, -1.2657e-01,
         -6.7472e-02, -1.4943e-01,  3.4114e-02, -5.5625e-02, -5.5094e-02,
          1.0176e-01,  1.2900e-01, -5.7207e-02,  1.8489e-02, -1.7177e-01,
         -7.2499e-02,  1.0768e-01, -8.6822e-03,  4.3501e-02, -1.1926e-01,
          1.1620e-01, -6.0562e-02,  7.4363e-02,  9.6805e-02,  2.6450e-02,
         -7.4517e-02, -6.7763e-02,  4.2590e-02,  9.4081e-02, -1.2800e-01,
          1.5388e-01, -7.2593e-02,  2.0515e-02, -7.4109e-02, -6.5941e-02,
          5.5008e-02, -1.8467e-02,  1.7082e-01, -2.2904e-02, -3.9810e-02,
         -7.6907e-02, -1.1589e-01,  1.8985e-02,  1.0085e-01, -4.1496e-02,
         -1.8363e-04,  9.5935e-02,  1.6373e-01,  1.7898e-01,  4.8950e-02,
         -4.9429e-02,  1.5055e-01,  1.2940e-01,  1.4366e-01,  1.1384e-02,
          2.9765e-03,  3.0897e-02,  1.1917e-01,  8.6979e-02,  4.1569e-02,
          8.4188e-03, -7.1886e-02,  1.1790e-01, -9.3509e-02,  8.5603e-02,
          7.8371e-03, -6.5506e-02,  6.0174e-02,  1.8929e-02, -1.6214e-02,
         -1.1463e-02,  1.1491e-01, -1.0321e-01, -1.6257e-02, -3.7207e-02,
          1.4291e-01,  1.2432e-01, -8.0419e-02,  4.0398e-02,  5.3929e-02,
         -1.1291e-02,  6.8221e-02, -9.7338e-02,  1.2540e-01,  5.1954e-04,
         -2.0926e-02, -7.1114e-02,  3.8985e-02,  4.7433e-02,  6.2325e-02,
         -8.1620e-02, -1.1341e-01, -5.2067e-02, -1.2000e-01, -1.2365e-01,
         -1.2876e-02,  6.0113e-02, -1.4734e-01, -1.0734e-01,  1.0377e-01,
         -4.3610e-02, -2.8074e-02, -7.4639e-02, -2.3198e-02, -1.0337e-01,
          6.1721e-02, -7.7622e-03, -1.3873e-02,  8.3889e-02,  1.1355e-01,
          5.4694e-02,  1.4811e-01,  1.6650e-01,  6.2975e-02,  2.4875e-02,
          1.1742e-03,  6.4305e-02, -1.0175e-01,  1.5465e-01, -1.5709e-01,
         -7.7609e-02,  7.2220e-02,  3.6013e-02,  6.5146e-02,  1.1933e-01,
         -2.6608e-02,  4.8176e-02, -1.3218e-01,  6.9404e-02,  4.2795e-02,
          2.7335e-02, -1.4227e-02,  2.9681e-02,  1.6850e-01, -7.7556e-02,
         -7.9868e-03,  8.7577e-02, -3.5371e-02, -4.9186e-03,  1.4551e-01,
          6.8346e-02,  7.0337e-02,  4.0058e-02,  1.3020e-01, -1.0048e-03,
          7.8430e-02, -5.9674e-02, -1.1097e-01, -1.2378e-03,  1.2719e-01,
         -8.9612e-02,  3.2255e-02, -2.3777e-02,  1.5967e-02,  8.6325e-02,
          1.0421e-01, -4.3836e-02, -5.4614e-02, -1.7539e-03,  1.1397e-02,
         -9.5316e-02,  8.0544e-02, -5.6412e-02,  2.2193e-02,  1.0408e-01,
         -1.2730e-01, -1.4134e-02, -8.3140e-02, -5.4082e-02,  1.0402e-01},
        '{ 1.0462e-01,  5.5912e-02,  2.2475e-02,  8.4921e-02, -1.4856e-01,
          5.8404e-02, -4.8843e-02, -1.9683e-01,  5.7130e-02,  6.0334e-02,
          9.2252e-02, -1.0334e-01, -9.0847e-02,  1.0375e-01,  9.5382e-02,
         -7.9893e-02, -2.8264e-03,  7.5851e-02, -2.1388e-02,  1.2075e-01,
          1.1494e-02, -5.6916e-03, -4.0958e-02, -1.0589e-01, -1.0480e-01,
          5.0822e-02, -7.8418e-02,  1.2484e-01,  1.8863e-02,  2.0842e-01,
         -1.2924e-01,  1.0633e-02,  1.2014e-01, -1.7110e-01, -1.3304e-01,
          4.0268e-02, -1.6550e-01,  3.9732e-02,  7.8918e-02, -6.8350e-02,
         -8.5062e-02,  1.3260e-01,  1.9768e-01, -5.3667e-02, -1.8484e-01,
          1.6657e-01,  1.8909e-01,  1.1502e-01, -6.2437e-02, -4.6191e-02,
         -1.4440e-01, -9.7840e-02,  4.9751e-02,  3.9487e-02,  6.5391e-02,
          1.0445e-01,  6.4356e-02,  1.1149e-01, -5.8553e-03, -1.2952e-01,
          9.2421e-02, -1.5047e-01, -1.5953e-01,  4.3969e-02,  9.3060e-03,
          9.7224e-02,  1.1137e-01,  9.8019e-02,  1.2295e-01,  1.3459e-01,
          9.2868e-02,  1.3642e-01,  3.4409e-02,  1.1821e-01,  2.4321e-02,
         -1.8108e-02, -1.2248e-02,  1.0898e-03,  9.3826e-02, -8.1069e-02,
          3.9522e-02,  9.1786e-02, -1.0026e-01, -1.1332e-01, -5.4090e-03,
         -4.5155e-02, -1.4195e-02,  8.7104e-03, -6.1931e-02, -1.9091e-01,
          8.4591e-02, -1.1129e-01,  4.4413e-02, -1.4524e-02, -7.5821e-02,
         -5.2530e-03,  2.9475e-02, -1.1881e-01,  8.5123e-02,  4.9304e-02,
          1.4664e-01,  6.9315e-02, -1.1166e-01, -6.6755e-02, -6.9803e-02,
         -3.1955e-02,  2.9478e-02,  8.0024e-02, -1.4012e-01, -1.6119e-01,
         -9.1033e-02,  1.5076e-01, -3.9324e-03, -3.6510e-02, -9.9332e-02,
         -6.8010e-02, -6.1545e-02, -5.8236e-02,  8.8007e-02,  6.4399e-02,
          1.1301e-01,  3.2695e-02,  3.8768e-02, -3.0055e-03,  1.6380e-02,
         -1.1562e-01, -2.4091e-02, -2.3264e-02,  9.4476e-03,  2.5565e-02,
          8.7966e-02, -6.2048e-02, -1.6759e-02,  2.9272e-02,  3.4806e-02,
          6.6357e-02, -1.9190e-02, -4.7540e-02, -8.3903e-02, -3.0007e-02,
          1.9689e-02, -3.0906e-02, -7.2460e-02,  6.0527e-02, -1.2488e-02,
          1.3124e-02, -3.2339e-02, -9.5436e-02,  1.1349e-01, -7.2709e-03,
          1.5660e-01, -6.8671e-02, -6.0996e-02, -6.8959e-03,  7.2012e-03,
         -3.6204e-02,  1.1481e-02, -7.2956e-02, -2.5415e-02, -1.8473e-02,
         -1.9012e-02,  1.1790e-01,  8.0304e-02, -7.8780e-02,  1.9455e-01,
         -1.5019e-01, -9.6611e-02, -1.0331e-01,  5.6559e-02, -5.2871e-02,
         -1.3073e-01,  9.3935e-02,  5.3328e-02,  1.2037e-01,  3.0520e-02,
          1.5313e-01, -5.1510e-02, -4.2098e-02,  1.3671e-01, -2.4334e-02,
          1.5802e-03, -8.7276e-02,  5.1891e-02,  2.6585e-02,  1.2165e-01,
          9.7108e-02, -4.3005e-03,  5.2800e-02,  9.6266e-02,  2.0401e-01,
         -1.4022e-01, -6.0818e-02,  3.5041e-02, -1.6783e-02,  1.9070e-01,
          4.6087e-03,  1.3249e-01, -1.4747e-01,  1.3294e-02, -6.7153e-02},
        '{-1.5222e-01, -6.7561e-02,  1.5426e-02,  9.6536e-02, -1.1951e-01,
          8.4443e-02, -1.8260e-03,  9.8736e-02,  1.2260e-02,  1.9015e-01,
          1.0834e-01,  9.7959e-02, -5.6845e-02,  2.0981e-02,  1.3232e-01,
          8.9747e-02, -4.7501e-02, -3.7362e-02,  9.2494e-02,  7.0258e-02,
          5.2028e-02, -1.4499e-02,  5.3633e-02,  5.4295e-02, -2.5867e-01,
         -1.5433e-01, -4.4588e-03, -1.0207e-01,  9.0710e-02,  2.5249e-01,
         -5.3175e-02,  1.7914e-01, -3.3909e-02,  1.8751e-01,  2.3133e-01,
         -6.9162e-02, -2.6095e-01, -7.9856e-02,  2.0416e-02,  1.1597e-01,
          1.9290e-02,  3.1099e-03, -1.0609e-01, -1.9615e-01, -4.5828e-02,
          6.6064e-02,  1.5913e-02, -1.1858e-01,  1.4307e-01, -9.3275e-02,
         -9.5062e-02, -2.7785e-02,  4.0832e-02, -3.6328e-02, -3.7492e-02,
         -4.8729e-02, -2.5628e-02, -1.0014e-01, -6.8503e-02,  1.3788e-01,
          3.0308e-02,  3.8600e-02, -2.8980e-02, -1.0579e-01,  1.0664e-01,
          3.1873e-02,  1.0204e-01, -8.8665e-02, -1.7527e-02,  1.6858e-01,
         -5.5927e-02,  1.2811e-01, -1.2347e-01, -1.4409e-02, -1.5197e-01,
          9.8755e-02,  3.0319e-02,  4.6364e-02,  2.6652e-02,  3.0654e-02,
          3.0754e-02, -1.0756e-01,  3.6842e-02, -1.3156e-01, -1.8758e-01,
          3.8657e-02,  7.7491e-03, -1.9623e-02, -8.0646e-02, -1.0141e-01,
         -2.5369e-02,  4.7559e-02,  1.0682e-02, -4.0776e-02,  5.4461e-02,
         -4.5845e-02,  1.2919e-01, -1.0957e-01,  6.0083e-02, -5.9299e-02,
          1.7969e-01,  7.8681e-03,  5.3093e-02,  3.6882e-03, -1.1798e-01,
          6.4874e-02,  7.3640e-02,  6.1603e-02,  1.0884e-01,  5.8016e-03,
         -9.9377e-02,  1.8146e-01, -3.7993e-02, -1.0274e-01,  1.0628e-01,
          9.1628e-02,  8.5800e-02,  9.7871e-02,  3.3126e-02,  3.0325e-02,
          1.0494e-01,  1.6686e-01,  1.1498e-02, -8.4864e-02,  6.6145e-02,
         -8.9542e-02, -1.9912e-02,  9.0930e-02,  1.8014e-01,  6.4940e-02,
          1.2240e-02,  5.8692e-02,  8.9378e-02,  2.0754e-01,  2.1850e-01,
          3.8890e-02, -6.5527e-02, -4.1840e-02, -6.1800e-02,  1.5751e-01,
         -2.0609e-02,  9.6067e-02, -4.1554e-03, -1.6190e-01, -1.0338e-01,
         -6.7240e-02, -4.2969e-02,  1.0534e-01, -9.8672e-02, -1.2384e-03,
         -8.7631e-02, -7.8457e-02,  6.5604e-02,  2.2271e-02,  1.0743e-01,
         -1.1978e-01,  1.1846e-01, -1.5884e-02,  1.2273e-01, -6.5392e-02,
          1.1162e-01, -1.0239e-01, -4.0727e-02, -1.3827e-01,  1.3463e-01,
         -3.2557e-02,  2.8214e-02,  7.5696e-02,  5.3907e-02, -5.4223e-03,
         -5.8512e-02, -4.0360e-02,  7.0368e-02,  6.6866e-02, -1.1528e-01,
          6.3396e-03,  1.3816e-01,  1.1698e-01, -1.1866e-01, -6.5179e-02,
          1.3375e-01,  1.6008e-01,  4.9569e-02, -1.0140e-02, -7.7426e-02,
          7.0863e-02, -2.4628e-02,  1.0117e-02, -2.0041e-02,  5.0042e-02,
         -3.1644e-02,  1.5590e-01, -1.0980e-01, -1.5786e-01,  9.8506e-02,
         -1.4182e-01, -4.9532e-02,  1.4506e-01, -8.5106e-02,  3.3883e-02},
        '{-5.0256e-02,  6.3192e-02,  1.9996e-01,  1.1655e-01,  1.1307e-01,
          1.1017e-01, -2.5312e-02,  8.5655e-02,  3.1730e-02,  8.9287e-02,
         -1.4118e-01, -3.3607e-02,  1.5853e-01,  1.4426e-01,  1.8070e-01,
          1.0072e-01,  3.0785e-02,  1.2124e-01,  3.0851e-02, -3.9615e-02,
          1.1781e-02,  2.1420e-02,  3.1121e-02,  4.9638e-03, -1.8167e-01,
         -1.0491e-02, -7.5721e-02,  4.2403e-02,  1.6411e-01,  1.0068e-01,
         -1.0722e-01, -4.1769e-02, -7.0649e-02,  3.3084e-02,  1.6875e-01,
          6.8855e-02,  6.9783e-02,  1.8452e-01, -3.2589e-02,  1.2855e-01,
          2.7707e-01,  1.5729e-01, -1.3746e-02,  1.1449e-01,  1.8423e-02,
         -3.8793e-02, -1.1698e-01, -1.9604e-01, -1.8722e-01, -1.5649e-01,
          3.6054e-02, -1.1058e-01,  3.4214e-02, -1.1757e-01, -1.1107e-01,
          1.3313e-01,  1.7057e-01, -1.3279e-01, -3.1795e-02, -1.4413e-02,
          7.1499e-02,  1.0499e-01, -2.0099e-03,  2.5961e-03, -1.1270e-02,
         -2.6850e-02, -4.8330e-02,  1.8913e-01,  2.2004e-01, -7.3375e-02,
         -7.7512e-02,  4.8522e-02,  1.4724e-01,  4.2599e-02, -4.2709e-02,
         -2.0643e-02, -8.3534e-02, -3.6779e-02, -2.2464e-01, -4.6108e-02,
          6.0895e-03,  1.1333e-01, -8.4593e-03, -2.3339e-01,  1.3991e-01,
          5.5417e-02,  5.6326e-03,  2.0142e-02, -6.0174e-02, -1.9973e-01,
          1.5335e-01, -9.0821e-02, -9.3370e-02,  2.0521e-01, -6.6878e-02,
         -6.8141e-02, -1.5545e-01, -3.6915e-02,  1.5245e-01,  1.6497e-01,
          1.3439e-01,  6.2486e-02,  9.0202e-02, -1.1143e-01,  4.9434e-02,
         -6.8721e-02,  1.9168e-01,  1.5553e-01, -6.5731e-02,  1.6067e-01,
         -8.4328e-02, -1.2561e-02,  4.8617e-02,  4.2411e-02,  7.8904e-02,
          1.0582e-01, -1.3064e-01, -9.1212e-02, -6.1116e-02, -1.2309e-01,
         -1.3172e-01, -4.4419e-02, -1.3811e-01,  6.0142e-02, -1.9665e-01,
         -7.0427e-02, -1.9547e-01, -3.4151e-02, -4.4074e-02, -3.4074e-02,
          3.7023e-02,  1.1027e-02,  6.0196e-02,  1.2392e-01,  6.1142e-02,
          1.3464e-01,  1.3035e-01,  2.1336e-01, -2.7834e-02,  9.1732e-02,
          1.9518e-01,  1.1082e-01,  1.0537e-01, -5.9180e-03,  7.9224e-02,
          8.9180e-03, -1.0968e-02, -2.8818e-02, -2.1608e-02, -4.4922e-02,
         -1.2696e-01,  9.4972e-02, -6.4793e-02, -5.5639e-02,  1.3226e-01,
          2.9846e-02, -1.1500e-02, -8.6793e-02,  4.2446e-02, -5.7696e-02,
         -1.2082e-01, -1.3443e-01, -9.9988e-02,  1.5300e-02,  6.4672e-02,
         -1.5195e-01, -3.5769e-02, -6.4963e-02,  6.2854e-02,  5.9694e-02,
         -1.1017e-01, -3.2999e-02,  1.3616e-01, -3.2208e-02,  2.0861e-02,
          1.7764e-01,  1.0178e-01, -3.1454e-02, -1.0605e-01,  1.1986e-01,
          2.0508e-02, -3.3899e-02,  3.9169e-02, -1.8933e-03,  1.8054e-01,
          1.4931e-01,  1.0155e-01,  2.9619e-02,  9.7362e-02,  1.7696e-01,
          5.4910e-02, -1.6746e-03,  6.9638e-02, -1.2575e-01,  9.0844e-02,
          1.1846e-01, -7.7898e-02, -3.1885e-02,  5.6247e-02, -1.9842e-02},
        '{-1.2456e-07, -4.0369e-23, -2.0633e-06, -3.1583e-06, -1.3525e-10,
         -1.2191e-06, -1.8002e-21, -2.8069e-06, -2.1943e-05, -2.4106e-05,
         -8.4760e-06, -1.6390e-05, -1.5577e-05, -1.3098e-05, -6.1570e-06,
         -8.0016e-06, -1.3463e-05,  1.0243e-05, -2.2868e-05, -2.7545e-05,
         -4.6277e-37, -1.1338e-10, -8.4102e-06,  8.9089e-22, -1.9637e-06,
         -5.0534e-07, -4.1027e-06, -7.9170e-07, -9.4795e-07, -1.4678e-06,
         -1.5419e-06, -1.1367e-07, -3.7681e-37,  2.5011e-08, -2.7670e-14,
         -1.7303e-07, -7.1106e-06, -1.6586e-17, -1.7031e-21, -8.9872e-06,
         -3.4040e-08, -6.1958e-11,  5.4264e-06,  9.2863e-22, -1.5716e-07,
         -1.3401e-05, -7.5327e-06, -1.6976e-05, -3.4927e-09, -1.5402e-06,
         -2.4853e-07, -6.3876e-10,  1.0066e-05, -4.3129e-06, -2.1984e-06,
         -1.3315e-12, -1.0426e-21, -1.2326e-05, -1.3728e-08, -2.6610e-21,
         -7.3503e-07, -3.6578e-06, -2.0768e-08, -1.8406e-05, -3.8993e-22,
         -7.8966e-06, -3.8401e-05, -1.2615e-05,  2.6139e-21, -3.1046e-07,
          4.1600e-21, -4.0875e-05, -2.5451e-06, -7.5374e-22, -8.9597e-22,
          1.4396e-37, -3.1975e-12, -2.2206e-05, -3.4751e-07, -7.6806e-15,
         -1.2140e-07, -4.8354e-06, -4.7727e-06, -3.5073e-09, -1.8510e-05,
          6.0507e-22, -1.2607e-07, -1.0381e-05, -2.1314e-05,  9.4235e-07,
         -1.7903e-05, -6.9285e-06,  6.2493e-06, -9.4118e-15,  1.1961e-06,
         -7.0292e-06, -1.7649e-07, -2.9062e-06,  6.4173e-10, -1.7383e-08,
         -1.5522e-08, -5.2622e-06, -3.5777e-12, -3.7765e-06, -9.7793e-09,
         -8.3732e-07, -3.6490e-06, -4.8500e-06, -1.1934e-05, -1.1411e-05,
         -4.5218e-06, -1.3711e-05, -1.5672e-05, -9.4318e-07, -1.6804e-05,
         -3.1114e-08, -2.0892e-21, -1.9808e-05, -1.0805e-05, -3.5075e-06,
         -1.3700e-05, -7.6793e-06, -1.0573e-07, -1.5158e-05, -1.9110e-05,
         -5.5744e-07, -1.6961e-07, -5.2763e-07, -2.8239e-06, -8.3657e-08,
         -1.4541e-08, -5.5828e-07, -4.3872e-30, -4.4126e-06,  2.3021e-21,
         -2.0620e-37, -5.0276e-06, -2.3314e-05, -8.2697e-06, -1.0443e-21,
         -8.5910e-06, -4.1628e-06,  1.1562e-22, -5.5960e-07,  1.5153e-05,
         -1.9880e-05, -2.0390e-05, -3.3008e-21, -3.8845e-07, -4.4346e-07,
          6.3957e-09, -3.6615e-06, -2.3344e-07, -5.4699e-07, -1.1395e-06,
         -3.0320e-11, -5.3596e-06, -1.7089e-05,  6.3707e-06, -7.5309e-13,
         -1.0547e-05, -9.3371e-06, -2.3835e-05, -2.6799e-05, -9.0807e-08,
         -7.4289e-06, -7.7055e-22, -1.8375e-05, -2.2443e-21, -1.7716e-05,
         -1.4447e-05, -2.5152e-05, -2.2044e-05, -1.4025e-05, -2.2625e-07,
         -1.1376e-09, -1.7190e-07, -3.1374e-12, -1.6383e-05, -2.1110e-05,
         -3.3910e-07, -2.7870e-06, -3.3566e-05, -2.6509e-06, -1.7148e-05,
         -2.2260e-05, -6.7880e-06, -2.8015e-05, -1.7970e-05, -2.0195e-05,
         -2.4483e-05, -1.9849e-05, -3.0580e-21, -2.6747e-21, -6.2903e-06,
         -1.4940e-05, -2.0499e-05, -4.9095e-06, -6.1622e-21, -4.6675e-06},
        '{-8.5956e-03,  1.6520e-01, -4.3676e-02, -6.0380e-02,  2.7198e-02,
         -1.4343e-01,  5.0575e-02, -3.6309e-02,  6.8852e-02,  1.1443e-03,
          1.4147e-01, -1.2944e-01,  8.4480e-02, -4.6224e-02,  1.1364e-01,
          4.6129e-03,  1.1266e-01, -6.1455e-02, -3.3296e-03,  1.0719e-01,
          9.8799e-02, -4.4840e-02,  2.4580e-01,  1.4822e-01, -6.0971e-02,
          1.2819e-02, -1.2013e-01, -9.0213e-02,  5.1802e-03,  1.1909e-01,
          9.8090e-03,  8.1329e-02, -7.7762e-03,  8.3111e-02,  2.6844e-02,
          1.0133e-01,  7.1508e-03,  7.8170e-02,  1.7027e-01,  2.2899e-01,
          1.6536e-02, -1.0610e-01,  3.3128e-02, -1.0044e-01, -1.1110e-01,
         -1.1933e-01, -1.0389e-02, -9.4053e-03, -1.4082e-01,  7.0381e-02,
          1.5656e-01,  1.2227e-01, -1.7628e-01, -1.5022e-01, -2.6298e-01,
         -1.2113e-01, -6.9477e-02, -1.0192e-01, -1.0044e-02, -4.3756e-02,
         -3.3352e-02, -5.9000e-02, -1.0310e-02,  2.0369e-02,  2.3517e-01,
          2.9882e-02,  1.1959e-01,  6.7571e-02,  1.0303e-01,  6.6379e-02,
         -1.3069e-01,  1.0354e-01, -5.9673e-02, -5.4007e-02, -1.0093e-01,
         -1.8240e-02, -8.4234e-03, -2.3412e-02, -9.4817e-02, -6.5893e-02,
         -1.3069e-01, -3.7199e-02, -1.0482e-01, -1.3382e-01,  2.5864e-02,
          2.6472e-02,  7.9097e-02, -7.9633e-03, -1.9736e-01, -5.9197e-02,
         -1.5063e-01,  2.0214e-01, -1.2911e-01,  1.1717e-02, -1.1798e-01,
          2.5745e-03,  1.2341e-01, -1.8588e-02, -3.1105e-02, -1.3069e-01,
          1.2728e-01,  7.8494e-02,  5.3728e-03,  5.2039e-02,  8.9327e-02,
          5.8980e-02,  1.5705e-01, -6.4626e-02,  3.9272e-02,  9.9686e-02,
          7.6254e-02,  1.6208e-01,  1.6889e-02,  5.7776e-02, -3.2104e-02,
          2.4450e-02,  6.5821e-02,  7.2017e-02,  3.8134e-02,  4.0975e-02,
          1.2684e-01, -2.5342e-02,  1.1154e-01,  8.3193e-02, -2.4769e-02,
         -9.9698e-02, -8.5550e-02,  3.6540e-02, -1.9420e-02, -1.4351e-01,
          1.4663e-01,  9.6775e-02,  1.0680e-01,  3.8173e-02,  2.2653e-01,
         -5.6228e-02, -6.6005e-02,  1.1594e-01,  9.2995e-02,  1.4191e-01,
         -5.4250e-02, -1.2948e-01, -6.7596e-02, -1.0192e-01,  9.1482e-02,
          1.1522e-01,  1.4685e-01,  8.4692e-02, -1.4575e-02,  4.8081e-02,
          1.2668e-01, -1.0020e-01,  1.7768e-01,  5.3500e-02, -8.0916e-02,
          1.0044e-01,  3.9665e-02, -4.1259e-02,  1.3827e-02, -5.5177e-02,
          7.2981e-02, -7.1671e-02, -1.4694e-01, -1.3026e-01, -4.4313e-02,
          9.8653e-02,  1.2815e-01, -1.3243e-02, -8.6468e-02,  1.9275e-01,
          1.1228e-01, -6.0126e-02,  4.7615e-02,  1.1700e-01,  2.5091e-02,
          3.4426e-02, -1.0540e-01, -1.0557e-03,  8.0394e-02,  2.8549e-02,
          1.5785e-01,  1.6847e-01, -1.3089e-02,  2.6370e-02,  2.2967e-02,
         -8.5866e-02, -5.7260e-02,  3.8421e-02, -1.9873e-01,  6.0403e-02,
          1.3456e-01,  4.6322e-02, -6.1827e-02, -1.5001e-01,  1.3874e-01,
         -1.3565e-01, -1.8256e-02,  1.0143e-01, -7.6609e-02,  1.1236e-01},
        '{ 2.9130e-02,  9.0895e-02, -3.7754e-02,  5.1117e-02, -1.1334e-02,
          2.3158e-02, -3.8385e-02, -8.8693e-02, -3.4608e-02, -9.3464e-02,
          9.6368e-02,  3.2819e-02,  1.0403e-01, -1.7005e-02, -4.5366e-02,
         -3.4744e-02, -4.2701e-02,  4.7034e-02, -9.8337e-03, -6.3887e-02,
          5.5524e-04,  5.6683e-03, -1.4857e-03, -1.3022e-02,  5.4332e-02,
         -2.7114e-02, -1.0581e-02,  3.2258e-02, -2.9637e-02,  2.2578e-02,
         -7.7047e-03, -2.3312e-03, -3.6279e-02, -1.1164e-02, -5.9790e-04,
         -4.8755e-06,  1.1285e-02,  1.0798e-02, -3.9189e-03,  2.6580e-05,
          4.8969e-02,  6.2495e-02, -6.6191e-03,  9.0235e-03, -8.6692e-03,
         -6.2750e-02,  2.2787e-02,  3.7403e-03,  2.9052e-02,  1.5597e-02,
         -1.4884e-02, -2.0096e-03,  1.7320e-03,  5.2476e-03, -3.3093e-02,
          4.4283e-03, -1.0550e-03, -2.8429e-03,  3.6443e-02, -2.7820e-02,
         -6.1070e-02, -3.2086e-03,  2.8216e-04, -4.1015e-02, -1.5337e-02,
          2.4851e-02, -3.6807e-02,  5.4319e-03,  2.4554e-02, -1.8462e-03,
         -1.4838e-02, -1.2738e-02, -7.4153e-03, -2.8484e-02, -3.6049e-02,
          1.8188e-03, -1.1903e-05, -3.2217e-04, -3.1369e-03,  3.8202e-03,
         -2.9923e-03, -2.1573e-05, -5.4782e-04, -4.1407e-03,  2.3906e-02,
         -3.4137e-03, -5.2670e-04, -1.5979e-03, -4.6409e-03,  9.8268e-04,
          9.6916e-03, -1.8519e-06, -2.2141e-04, -3.2061e-03, -1.6046e-03,
         -4.1565e-04, -1.0120e-04, -4.7775e-04,  1.9264e-02, -1.7115e-03,
          8.3612e-04, -5.6706e-02,  2.1603e-03, -6.0862e-02,  6.6923e-02,
         -6.0350e-02,  9.1895e-02,  1.7565e-02,  3.9560e-02,  2.4128e-02,
          1.0016e-01,  2.3453e-02, -9.6182e-02, -4.3017e-02, -9.9125e-02,
          9.2874e-02, -4.5605e-02, -1.1683e-01,  6.2154e-02,  9.4725e-02,
         -2.4413e-02, -2.5439e-02, -2.7337e-02, -9.3780e-02, -3.4397e-02,
         -6.1727e-05, -2.2494e-05, -2.4622e-04, -7.9220e-04,  1.2988e-03,
          1.4439e-02, -5.2874e-03, -1.2896e-03, -6.8286e-03,  2.6041e-02,
         -5.9324e-02,  3.2874e-02, -8.6153e-03, -2.2723e-03, -3.2964e-02,
          4.7426e-02,  6.9700e-02, -6.4146e-03, -4.8547e-02,  7.1853e-03,
          1.5664e-02,  1.1253e-03,  9.4419e-03, -2.6161e-02, -1.8787e-02,
         -3.8552e-03, -6.8933e-02, -1.8803e-02, -4.5149e-02,  3.4997e-03,
          1.5789e-02, -1.8201e-02,  9.9902e-03, -2.7449e-02,  2.4407e-02,
         -7.8567e-02, -8.1569e-02, -6.1630e-02,  4.4235e-02, -5.0129e-04,
         -3.5589e-02,  6.7468e-02,  8.2058e-02, -6.2084e-02,  4.7012e-02,
         -1.9977e-03, -9.4358e-04, -1.7262e-03,  1.9442e-02,  1.0612e-02,
         -1.4766e-02,  6.0438e-02, -6.6456e-03,  2.8507e-02, -9.1126e-02,
         -2.5263e-02, -1.0390e-01,  7.5936e-02,  2.6491e-02,  7.1702e-03,
          9.2926e-02,  8.1045e-03,  3.4936e-02, -9.9765e-02, -7.1448e-02,
          2.4563e-02,  2.5627e-02,  3.7730e-02, -6.3243e-02, -4.3298e-03,
         -1.3072e-02, -4.1725e-02,  1.4723e-02, -2.9520e-02,  9.5070e-04},
        '{-1.3111e-01, -2.7134e-02, -5.3969e-02, -1.2351e-01, -5.5260e-02,
          2.1546e-02, -1.0341e-01, -5.6272e-02,  2.2278e-04,  1.9161e-01,
         -2.4615e-02, -9.4086e-02, -6.0662e-02, -1.3698e-01,  1.2766e-01,
         -1.3351e-01,  1.3106e-01,  5.5249e-02,  5.5630e-02,  1.7890e-01,
         -2.9327e-02, -1.3915e-01,  2.4433e-01,  1.3673e-01,  1.4828e-02,
         -1.3373e-01, -1.4525e-01,  8.6193e-03, -2.3880e-02,  5.2312e-02,
         -2.1413e-01, -7.7618e-02, -2.4060e-01,  9.4499e-02,  7.9261e-02,
         -1.2028e-01, -2.2705e-01, -1.7078e-01,  2.9228e-02,  8.5104e-02,
          2.4512e-02, -2.8576e-01, -2.4430e-02, -1.4974e-01,  7.2398e-02,
         -7.8909e-02, -2.1532e-01, -2.1774e-01, -1.2415e-01, -3.6348e-02,
         -8.5747e-02,  3.7116e-02, -1.1186e-01,  2.9327e-02,  7.8370e-02,
          1.4604e-01, -2.6460e-02, -1.6506e-01, -1.6354e-01,  2.9152e-02,
         -1.0064e-01,  8.6690e-02, -8.3970e-02, -6.6330e-02,  1.3288e-01,
         -3.8421e-02,  6.6606e-02, -2.5783e-02, -7.4236e-02, -6.3454e-02,
          9.5953e-02,  2.0227e-03, -2.4566e-02, -1.6798e-01, -8.5606e-02,
         -4.9725e-02,  1.1042e-01, -3.8817e-02, -3.0128e-02,  1.1265e-01,
         -9.4557e-02,  1.2571e-01, -8.6222e-02, -8.9427e-02,  5.9358e-02,
          3.6900e-03,  1.6202e-01, -2.8019e-02,  4.4849e-02, -1.0218e-02,
          3.8027e-02,  1.2694e-01,  2.5736e-02, -3.7569e-02,  5.7899e-02,
          1.0797e-01,  1.1213e-01, -2.4379e-02, -3.7687e-02, -3.9912e-04,
         -2.2572e-02,  7.1400e-02,  1.0421e-01,  1.2115e-01,  1.5492e-01,
         -5.6311e-03,  7.0808e-02,  4.3777e-02, -9.1709e-02,  9.6312e-03,
          1.2733e-01,  1.6340e-01,  8.0315e-02,  2.0420e-02,  1.8679e-01,
          3.3149e-02,  8.1568e-02, -7.8436e-03, -6.6470e-02,  4.5042e-02,
          2.1867e-02, -4.5204e-02,  5.4740e-02,  1.4830e-01,  1.4443e-01,
          9.8896e-02, -1.1690e-01, -5.1766e-02,  6.6678e-03,  2.1325e-01,
         -9.2724e-02, -4.0062e-02, -2.0216e-01, -1.6257e-02,  3.3434e-02,
          3.1319e-02,  1.2021e-01,  7.3752e-02, -6.7759e-02,  1.7746e-01,
          2.6692e-02, -5.8696e-02, -1.1438e-01, -1.6999e-01,  7.2777e-02,
         -8.9150e-02, -6.0807e-02,  4.0129e-02,  1.2149e-01,  1.1508e-01,
          5.6107e-03, -1.3867e-03,  1.3226e-01,  6.8535e-02, -5.4502e-02,
         -4.8740e-02,  1.6363e-01,  7.2184e-02,  1.1037e-01, -7.4951e-02,
         -7.0401e-02, -2.9094e-02,  1.1275e-01, -6.3704e-02, -5.3379e-02,
          1.3250e-01,  1.5186e-01,  5.6940e-02,  2.5846e-02, -8.0392e-02,
          2.0852e-02,  5.3642e-02, -2.6699e-03,  1.2060e-01,  7.9969e-03,
          2.4330e-02,  3.7631e-02, -3.7829e-04,  5.5362e-02, -7.4001e-02,
          8.3330e-03,  1.4949e-01,  1.2838e-02, -9.1993e-02, -2.3398e-02,
          8.4325e-02, -3.7318e-02,  7.5846e-03, -1.6531e-01, -2.6435e-02,
          3.7596e-02,  3.5381e-04, -5.9586e-02, -1.0254e-01, -7.4183e-02,
          5.7044e-02,  4.7785e-02, -5.2284e-02, -3.3539e-02, -1.2723e-01},
        '{ 1.1498e-02,  6.4130e-02, -3.3209e-02, -6.2997e-02, -8.0101e-02,
          7.7619e-02,  1.0265e-01, -8.1776e-02,  5.1295e-03,  7.3879e-03,
          5.8348e-02, -3.8196e-02,  7.6243e-02, -5.0677e-02, -1.1313e-01,
          1.4756e-01, -3.5050e-02,  6.1323e-02,  4.9891e-02,  3.2955e-04,
         -5.0375e-02,  9.8099e-03,  3.0623e-02, -1.3894e-01,  1.0491e-01,
         -5.7061e-02,  2.1900e-01,  3.0119e-02, -2.0857e-01, -2.9143e-01,
          2.5150e-01,  1.6883e-01,  4.1055e-02, -1.7398e-01, -3.3109e-01,
          2.9431e-02,  2.8254e-01,  1.5930e-02, -7.0172e-02,  5.3031e-02,
         -9.3666e-02,  2.7497e-01,  1.4677e-01,  1.0235e-01,  6.1203e-02,
          1.8502e-01,  9.8089e-02,  9.9705e-02,  1.0342e-01, -6.5770e-02,
         -6.3175e-02, -1.5163e-01, -4.2291e-02,  2.1397e-01, -3.4487e-02,
          8.1549e-02, -3.5922e-02,  3.0908e-02,  5.3494e-02, -1.4619e-02,
          6.0430e-02,  7.9218e-02,  1.1676e-01,  8.2306e-02, -5.9488e-02,
         -1.4737e-01,  8.6757e-02,  1.9215e-01, -8.4287e-02,  5.8290e-02,
          3.3623e-02,  2.3479e-02,  2.9407e-03, -5.3874e-02,  1.2804e-02,
         -6.4322e-04,  1.8929e-02, -1.4850e-02, -1.3265e-01, -1.7522e-01,
         -1.3212e-01, -8.1572e-02, -9.6765e-02,  6.9295e-02,  4.6555e-02,
         -4.9046e-02, -6.2568e-02, -1.6729e-01,  1.8012e-01, -3.7611e-02,
          3.2044e-02,  2.1058e-02,  3.6116e-02, -2.1866e-02,  8.5918e-03,
         -7.0945e-02,  3.4605e-02,  1.4359e-01, -1.0955e-01, -9.2415e-02,
          1.1784e-01,  9.6042e-02,  1.2684e-01, -6.8643e-02, -4.7040e-02,
          1.0797e-02,  9.5076e-02, -7.4478e-02,  1.2531e-01,  1.0057e-01,
         -6.9028e-03,  3.1550e-02, -1.6234e-02,  6.6395e-02,  1.2982e-01,
         -1.1941e-01, -8.9694e-02, -3.8328e-02,  5.8557e-02,  1.4191e-03,
          3.0061e-02, -4.0378e-03, -4.9661e-02,  4.0404e-02, -1.3534e-02,
         -7.0091e-02,  6.6305e-02, -2.8463e-02,  1.0868e-01, -1.1468e-01,
          1.8444e-01,  1.1864e-01,  9.3278e-02,  2.0721e-02, -2.2837e-01,
          1.4050e-03,  4.1564e-02,  1.2040e-01, -1.3386e-01, -1.7181e-01,
         -1.0751e-01,  7.6685e-03,  2.3262e-01,  5.9588e-02,  1.3815e-01,
          1.0138e-01, -3.6256e-02,  1.3181e-02, -1.0070e-01,  7.0614e-02,
         -6.8003e-02,  6.5035e-02,  4.5719e-02, -2.2909e-02,  6.9223e-02,
          6.2248e-02, -1.6170e-02,  9.4112e-02,  1.8800e-01, -7.3584e-02,
         -1.2957e-01,  5.9598e-03,  1.6713e-01, -1.2769e-03,  1.5785e-01,
          2.8021e-03,  6.3614e-02, -6.1177e-02, -5.7434e-02,  5.9365e-02,
          8.3132e-02, -9.4175e-02,  2.1573e-02, -2.0312e-02,  3.1536e-02,
          1.7236e-02,  8.7783e-02, -1.0284e-01, -8.3313e-02, -1.3172e-02,
          3.2336e-02,  1.3747e-01, -3.1593e-02,  1.0538e-01, -2.0358e-02,
         -5.2410e-02,  9.0767e-02,  5.0979e-02, -1.9826e-02, -7.8530e-02,
         -4.7504e-02, -8.5999e-02, -1.2984e-02,  5.4173e-02, -7.8622e-02,
          1.2479e-01,  1.2671e-02, -1.4875e-01, -3.5039e-02,  1.3335e-01},
        '{ 1.1961e-01,  6.7360e-02,  5.9692e-02,  2.3813e-01,  1.1161e-01,
          1.7080e-01,  1.5014e-01,  2.1560e-01,  2.2540e-01,  4.7562e-02,
         -3.7640e-02, -3.7536e-02, -1.6107e-01,  3.8185e-02,  3.1127e-02,
         -1.5869e-01,  1.9637e-01,  1.0718e-01, -1.2350e-01, -9.2820e-02,
         -7.1038e-03, -1.3680e-01,  9.2024e-02, -1.7923e-01, -1.1015e-01,
          9.8425e-02,  1.1131e-01, -1.6956e-02, -8.0357e-02,  4.1242e-03,
          7.4095e-02,  1.4972e-02,  2.1502e-01,  9.4765e-02, -2.0937e-01,
         -8.3794e-02, -1.6949e-02,  6.9073e-02,  6.1410e-02, -1.0539e-01,
         -1.8808e-01, -1.5903e-01,  8.3933e-02, -1.6387e-01,  1.6365e-02,
          8.6764e-03,  7.5510e-02, -1.2473e-01,  1.0658e-01,  1.7296e-01,
         -1.5695e-01, -2.9442e-02, -1.8041e-01, -1.5469e-01, -1.4519e-01,
          1.2953e-02, -6.1090e-02,  9.9326e-03, -1.9114e-02,  1.0391e-01,
          1.0348e-01, -1.4325e-01,  8.2214e-02,  1.6981e-01,  2.3483e-01,
          7.2589e-02,  1.2146e-01, -1.9417e-01,  7.3989e-02, -4.3222e-02,
         -9.8424e-02, -1.9788e-02, -1.0855e-01, -2.1877e-02, -2.1910e-02,
         -6.4820e-02, -9.1353e-02,  4.8416e-02, -1.2789e-01, -2.2592e-01,
         -1.4145e-01, -7.2042e-02, -5.7844e-02, -1.3440e-01, -1.8757e-01,
          3.0859e-02,  3.7334e-02,  1.3541e-01, -6.4771e-02,  1.0614e-01,
          2.4365e-02,  2.1177e-02, -1.6551e-02,  2.1257e-02,  1.2052e-01,
         -1.5703e-02,  9.6600e-02,  4.3599e-02, -4.3730e-02, -1.2643e-01,
          8.7158e-02,  1.3021e-01, -3.9914e-02,  2.6050e-02, -1.0471e-02,
          1.2814e-01,  1.5271e-01,  1.5382e-01,  3.3318e-02,  6.8839e-02,
         -7.7395e-02,  1.1369e-01,  5.6439e-02, -3.4175e-02,  1.2901e-01,
         -1.1987e-01,  3.4505e-02, -1.7753e-02, -1.4207e-01,  1.1986e-01,
          6.7088e-02, -1.7945e-02,  3.9763e-02,  5.7131e-02,  4.8395e-02,
         -7.8767e-02, -7.8488e-02, -1.2824e-01, -7.5568e-02, -6.4027e-02,
         -1.0463e-01, -5.5223e-02, -1.8471e-02,  5.2783e-02,  9.2817e-02,
          8.6295e-03, -2.4290e-02, -1.0398e-01, -3.1405e-02,  9.1889e-02,
         -8.5390e-02,  2.8128e-02, -1.4198e-01, -7.4131e-02,  3.7135e-02,
         -1.4127e-01, -1.0273e-01, -4.9306e-02,  4.6190e-02, -1.1542e-01,
         -4.4237e-02,  1.1752e-01,  1.3413e-01, -3.7721e-02, -4.8942e-02,
         -6.2890e-02,  6.7340e-02,  3.0560e-02,  2.0848e-01, -5.8462e-02,
         -7.7328e-02,  1.2088e-02, -1.6234e-01,  6.5093e-02,  8.5387e-02,
          1.4439e-01,  1.2601e-01, -1.0174e-01, -1.1775e-01, -8.7240e-02,
         -1.4889e-01, -1.0350e-01, -7.9075e-02,  1.3463e-01, -1.9976e-01,
         -1.5999e-01,  8.2629e-02, -6.0677e-02,  1.0670e-01,  1.2539e-01,
          1.1312e-01,  1.5970e-01,  1.2315e-01,  7.2279e-02,  1.9915e-01,
          1.0402e-01, -9.8690e-02, -3.7119e-02, -4.7131e-04,  2.0556e-01,
         -2.2398e-02, -9.9080e-02, -7.3436e-02,  8.2252e-03,  4.7946e-02,
          1.1992e-01, -6.0111e-02, -4.2898e-02,  4.1206e-02, -1.6270e-01}}
;

real fc1_bias_re[64] = 
      '{-1.6529e-02,  4.6535e-03,  1.4074e-02,  4.8890e-02,  2.7984e-02,
         3.7829e-02,  3.0358e-02,  3.4421e-03,  2.4707e-02,  5.4348e-03,
         2.6795e-05,  2.8556e-03,  1.9299e-02,  4.9210e-02,  1.8319e-02,
        -8.9894e-03, -1.4062e-02,  1.9371e-02, -4.2791e-03,  1.9258e-02,
        -2.2905e-02,  1.6871e-02,  1.2313e-02,  1.3832e-02, -1.4009e-02,
         1.3131e-02,  2.2812e-02,  4.9683e-03,  4.1242e-02,  2.5681e-03,
         2.0147e-03, -1.9226e-03, -3.8133e-03, -8.6936e-03,  1.2835e-02,
         2.2934e-02,  1.1112e-02,  1.6311e-02, -2.7403e-02, -1.5499e-02,
        -2.1783e-03,  5.4207e-04,  5.7142e-03,  3.5094e-02, -2.9501e-03,
         2.1615e-02,  1.3742e-02, -6.1479e-03, -2.0175e-02,  4.5612e-03,
         7.7907e-03,  3.6275e-03, -1.0665e-02, -4.0339e-03, -1.5490e-02,
        -1.8666e-02, -4.7386e-03,  9.6818e-03,  2.2946e-21,  1.1161e-02,
         1.1104e-03,  1.0647e-02, -4.5903e-03,  6.4241e-03};

real fc2_weights_re[10][64] = 
     '{'{ 1.5505e-01, -2.9713e-02,  1.3664e-01, -2.3565e-01, -9.1041e-02,
          9.4507e-02,  2.9844e-01,  2.6090e-01, -3.7817e-01,  2.1072e-01,
          3.0684e-03, -7.6007e-02, -1.9224e-01, -2.1731e-01,  1.8155e-02,
         -6.6715e-02, -7.3174e-02,  4.2511e-02,  2.0613e-01, -3.0824e-01,
         -9.4993e-03,  6.6291e-02, -5.8045e-03, -1.0618e-01,  1.6842e-01,
          8.0115e-02, -2.0660e-02,  1.0884e-01,  1.1105e-01,  9.6579e-02,
          2.3574e-01,  1.1921e-01,  7.9128e-02, -2.2683e-02,  2.3366e-01,
         -2.8015e-01,  1.2433e-01, -3.5657e-01, -3.5707e-01,  3.7041e-01,
          4.9643e-02,  3.6617e-02,  1.7980e-02, -1.4375e-01, -5.3712e-07,
          1.7816e-01, -3.4215e-01,  2.9401e-01,  1.2915e-01,  6.2508e-02,
         -6.8198e-02, -1.1531e-01, -8.1898e-02,  2.9580e-04, -2.5636e-01,
         -1.5987e-01,  2.8674e-01, -5.4382e-02,  4.9768e-06,  2.4235e-01,
          2.2498e-04,  2.2157e-01, -2.8057e-01,  2.6698e-01},
        '{-3.3480e-01, -3.4808e-01, -1.4608e-01,  3.1609e-01, -7.1175e-03,
          1.6684e-01,  7.4646e-02, -3.2223e-01, -8.4993e-02,  3.7568e-01,
          6.2197e-03,  2.3722e-01,  2.3181e-01,  1.4315e-01, -3.1695e-02,
          4.4405e-02, -1.6535e-01,  8.9789e-02, -3.7132e-01, -1.0544e-01,
         -2.6494e-01, -2.1924e-01,  2.0656e-02,  1.9498e-01, -2.4235e-01,
         -3.0584e-01,  2.2181e-01,  1.2359e-01, -1.3884e-01, -1.8952e-01,
         -7.3897e-02, -2.0815e-04,  2.0781e-01,  1.9462e-01,  2.1778e-02,
          5.3716e-04, -2.0005e-01,  6.2935e-02, -1.3402e-01, -2.4542e-01,
         -9.2537e-05, -2.3338e-02, -3.7370e-01,  2.7430e-01, -4.5061e-04,
         -7.2898e-02, -1.8775e-01, -9.3686e-02,  5.1293e-02,  1.6841e-01,
          7.8830e-02,  7.1826e-02,  1.9306e-01, -1.4471e-03,  1.0724e-02,
         -2.6640e-01, -3.9159e-01, -2.3422e-01, -5.5269e-10, -3.5688e-01,
         -5.5385e-07, -3.3119e-01, -1.1121e-01, -2.9971e-01},
        '{ 3.2743e-01,  2.5521e-01, -2.9408e-01, -1.0120e-01, -4.3992e-01,
         -1.7650e-01,  2.8207e-01, -6.5359e-03, -1.6879e-02,  1.6515e-01,
          2.2009e-03, -6.3591e-02, -1.3845e-01,  2.2096e-02, -2.9218e-01,
         -3.5285e-03, -3.0368e-01,  2.5802e-01, -1.5643e-01,  2.3268e-02,
         -1.5694e-01, -1.3185e-01, -1.7019e-01,  1.9468e-01, -1.7092e-01,
          1.5519e-01, -1.0203e-01,  3.1554e-01, -3.4307e-02,  3.2629e-01,
         -5.7628e-02, -7.3535e-03,  1.9810e-01,  6.3925e-02,  1.7914e-01,
         -2.9108e-01, -8.9571e-02,  1.9791e-01, -2.7942e-01, -2.4743e-01,
          5.2378e-03, -3.5351e-01,  2.1471e-01, -2.4713e-02, -4.5803e-04,
         -1.1556e-01,  1.4331e-01, -8.7567e-02, -2.2878e-01,  7.4509e-02,
         -1.8287e-02,  2.9757e-01,  1.1834e-01, -1.0764e-02, -2.8249e-01,
         -1.7843e-01, -1.1308e-01, -2.9518e-01, -3.1211e-04, -5.7219e-02,
          1.7444e-04, -1.4064e-01,  1.8742e-01, -1.1341e-01},
        '{ 1.2712e-01, -1.1703e-01,  8.8066e-02, -1.3318e-01,  1.6133e-01,
          4.3562e-02, -8.0526e-02, -2.6987e-02,  3.5309e-02,  9.4382e-02,
         -1.1693e-02, -2.5140e-01, -2.9891e-01, -2.4777e-01,  2.8159e-01,
          2.9000e-01, -4.8158e-02, -8.7344e-02, -5.8539e-02, -1.0062e-01,
          3.8375e-01, -3.9222e-01,  1.2375e-02, -1.7225e-01,  1.0132e-01,
          4.1097e-02,  9.6104e-02, -3.0193e-01, -1.3294e-01, -1.4117e-01,
         -2.0309e-01, -9.7932e-04,  5.3322e-02,  7.3612e-02, -3.1055e-01,
         -1.4376e-01, -1.6367e-01,  2.9125e-03,  2.5278e-01,  1.0431e-01,
         -5.1162e-03, -6.5047e-02, -7.8562e-02,  7.8070e-04, -6.8838e-03,
          7.6836e-02, -4.5850e-02,  2.9072e-01,  2.3198e-01,  2.0537e-01,
         -1.2303e-01,  1.2775e-01,  1.4183e-01, -8.5445e-03,  9.2802e-02,
          2.1829e-01,  1.0329e-01,  1.1455e-01, -4.2605e-07, -4.2228e-02,
         -7.0082e-04, -2.6023e-01,  1.2706e-01,  1.0188e-01},
        '{-7.3402e-02,  2.8730e-01, -2.3309e-01, -1.6068e-01, -1.6860e-01,
          1.3800e-01, -3.9337e-01,  3.0914e-01,  2.2398e-01, -5.5053e-02,
         -1.2055e-02,  2.0579e-01,  3.0542e-01, -1.0168e-01, -3.8288e-01,
         -1.0612e-01,  3.2951e-01, -3.6486e-02,  2.4816e-01, -2.5836e-01,
         -4.2178e-01,  2.3298e-01, -2.9986e-01, -3.2511e-01,  2.6415e-01,
          1.1415e-01, -2.7283e-01, -1.5238e-01,  2.3819e-02,  2.9310e-02,
         -4.3723e-02, -2.5599e-02,  1.8989e-01,  3.3380e-01, -2.1717e-01,
         -2.2847e-01,  2.2157e-01, -1.6190e-01,  1.1043e-01, -4.9838e-02,
         -4.7444e-03, -4.8071e-01, -3.0461e-01,  8.4906e-02,  4.7424e-03,
          9.4778e-02, -2.9328e-01, -2.6714e-01, -2.1956e-01,  1.1374e-01,
         -8.6819e-05, -3.4391e-01, -4.9426e-02,  3.2632e-03,  2.8001e-01,
          4.6057e-02, -1.9558e-01,  2.0122e-01, -2.8156e-08, -2.1715e-01,
         -8.9768e-02, -2.3179e-03,  1.0534e-01, -3.7509e-01},
        '{-6.1658e-02,  3.9622e-02,  8.7758e-02,  2.5282e-01,  2.6209e-01,
          2.9238e-01,  8.8519e-02,  2.1992e-01,  5.2253e-02, -2.9094e-01,
         -7.8857e-02,  2.3538e-01, -2.6965e-02,  8.9596e-02,  2.6082e-01,
         -5.4927e-02, -2.5189e-01,  1.0762e-01, -8.1056e-02, -3.3449e-01,
         -1.4700e-01,  7.1715e-02,  8.0757e-02, -2.4162e-01, -1.2631e-01,
          1.1022e-01,  1.7477e-01, -2.7211e-01,  2.9908e-01, -1.6236e-01,
         -3.7937e-01,  2.6637e-03, -1.0208e-01, -1.7840e-01, -2.0066e-01,
         -7.0357e-03,  2.6208e-01, -1.7005e-01, -2.6578e-02, -1.8724e-01,
          5.2663e-02, -2.0845e-01, -1.5116e-01, -9.0430e-02,  6.5000e-05,
          1.1956e-01,  8.9190e-02,  1.0830e-01, -2.0956e-01,  8.3619e-02,
         -3.4131e-02, -2.0637e-02, -3.6615e-01, -7.7294e-03, -2.4500e-01,
         -6.0345e-02,  1.7270e-01,  3.0262e-01, -4.8847e-05,  1.0729e-01,
         -4.0827e-05, -3.1912e-03, -1.9434e-01, -2.2204e-01},
        '{-5.5123e-02, -2.9486e-01,  1.4136e-01,  2.3271e-01, -1.7263e-01,
         -3.4535e-01,  2.0630e-01,  2.9239e-01, -5.4343e-02, -1.7847e-01,
         -1.2994e-02, -1.1856e-01,  1.6782e-01, -7.7894e-02,  1.0552e-01,
         -2.9074e-01,  2.0560e-01,  3.3414e-01, -1.5032e-01, -2.6081e-01,
         -1.4861e-01, -8.0899e-03, -5.0503e-02, -3.7214e-01, -2.2346e-01,
          4.9910e-02,  2.7343e-01, -1.9126e-01,  2.4268e-01, -3.0246e-01,
          1.1586e-01, -9.9376e-04, -3.2446e-01,  1.8355e-02,  2.7994e-01,
         -8.2582e-02,  2.6460e-03,  5.8563e-02,  1.1648e-01,  2.6693e-01,
          1.2307e-04, -2.6189e-01, -3.2682e-01, -1.1633e-01,  9.3236e-06,
         -4.3249e-01,  8.9325e-02,  1.8136e-01, -7.5197e-03,  1.1873e-01,
         -4.0054e-01, -3.4182e-01,  3.0652e-01, -2.9905e-03,  2.4079e-01,
          1.8192e-01,  3.2774e-01, -1.6242e-01,  5.7795e-03, -7.1860e-02,
          3.5319e-05,  1.3920e-01, -2.6431e-01,  1.4709e-01},
        '{-2.0760e-01,  7.3112e-02, -1.0314e-02,  1.4074e-01, -7.2170e-02,
          1.1377e-01,  1.3416e-01, -2.6590e-02,  9.2885e-02,  2.8403e-01,
          1.4794e-02, -1.3603e-01,  2.5975e-01, -3.0335e-01,  3.1689e-01,
         -3.5107e-01, -6.9212e-04, -3.1493e-01, -1.9759e-01,  2.6161e-01,
         -3.2760e-01, -2.5175e-01,  1.3964e-01,  2.7885e-01,  8.7769e-02,
         -3.0889e-01, -3.7567e-01, -1.5118e-01,  1.4369e-02,  2.4523e-01,
          5.3049e-03, -2.2966e-01, -2.7172e-01, -6.1106e-02,  1.0286e-01,
         -4.0451e-01,  7.3992e-02,  8.1419e-02, -1.7416e-01,  1.2923e-02,
          9.7200e-10,  6.2738e-02,  3.2858e-01,  1.3796e-01, -4.8537e-02,
          2.3933e-01, -2.4657e-01, -1.8340e-01,  7.8541e-02,  2.4573e-01,
          1.7968e-01,  1.9339e-01, -1.2152e-01, -3.1217e-02, -1.1169e-01,
         -1.5854e-01,  9.1594e-02,  2.7946e-01, -1.6261e-03,  2.6385e-02,
          9.6035e-03, -4.2581e-02,  1.8248e-03,  3.3531e-01},
        '{ 2.5627e-01,  1.5938e-01, -2.5920e-01, -6.0286e-02, -2.9377e-01,
         -5.8784e-02,  1.1950e-01, -1.2017e-01, -1.8935e-01,  1.4765e-01,
         -6.0156e-02, -1.2878e-01,  2.5058e-01,  1.6398e-01, -2.8477e-01,
          1.9260e-01,  1.6867e-01, -5.6877e-02, -1.2058e-01,  7.3404e-02,
          6.0162e-02, -5.4070e-02, -6.0996e-02,  1.9520e-01,  2.2993e-01,
         -2.7253e-01,  2.8456e-01,  2.8420e-01, -3.5255e-01, -2.6227e-01,
          1.1489e-01, -2.5000e-03, -3.2588e-01,  2.6284e-01, -3.2800e-01,
          5.0247e-03,  4.9309e-02, -6.8976e-02,  1.4313e-01, -1.0028e-01,
          1.1007e-04,  1.7410e-01, -7.8866e-02, -2.0960e-01, -3.1314e-03,
         -2.8536e-01, -7.5696e-02, -3.5490e-01, -3.4097e-01, -3.6887e-01,
         -1.3042e-02,  3.3459e-02,  2.0021e-01,  1.8349e-02, -1.8870e-01,
         -2.1352e-01, -5.2145e-02,  3.1462e-01, -8.4617e-04,  1.0036e-01,
         -4.2114e-03,  1.0722e-01, -6.4816e-02,  5.4949e-02},
        '{ 1.2920e-01,  2.0818e-01, -3.8263e-01,  3.1584e-01,  2.2736e-01,
          2.6812e-01, -3.6159e-02, -4.2398e-02,  1.6969e-01, -4.0180e-02,
         -5.8909e-03, -4.3318e-03, -1.1733e-01, -7.2175e-02, -3.0151e-01,
         -2.8546e-01,  9.5526e-02, -3.9331e-01,  1.4224e-01,  2.7859e-01,
         -9.8346e-02, -1.2108e-01,  3.3258e-02, -1.0942e-01, -7.1416e-02,
          2.7228e-01, -1.6748e-01,  7.2192e-02, -1.0903e-01, -3.3570e-02,
          3.1694e-01, -1.1001e-02, -1.2975e-01, -2.2294e-01, -9.7771e-02,
          1.8116e-01, -9.7278e-02, -1.8572e-01, -1.5879e-01,  5.7298e-02,
         -6.2813e-05, -3.2273e-01, -6.7278e-02,  1.2552e-01, -4.6552e-04,
          2.4132e-01,  1.4291e-01, -1.8976e-01, -7.3817e-02, -2.7829e-01,
         -3.3398e-01, -2.9183e-01,  2.3535e-01, -1.9732e-02,  2.2260e-01,
          1.0663e-01, -1.4513e-01,  1.4706e-01,  9.3050e-04, -2.7357e-01,
          5.7909e-03, -4.2781e-01,  1.1080e-01,  2.9883e-01}};

real fc2_bias_re[10] = '{-0.0282,  0.0321,  0.0077, -0.0252, -0.0009,  0.0377, -0.0116, -0.0033, -0.0133, -0.0028};


